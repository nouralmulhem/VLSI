
// 	Thu Dec 22 23:04:39 2022
//	vlsi
//	localhost.localdomain

module Register__parameterized0 (clk_CTSPP_21, clk_CTSPP_62, clk_CTSPP_72, in, clk, 
    out);

output [63:0] out;
input clk;
input [63:0] in;
input clk_CTSPP_21;
input clk_CTSPP_62;
input clk_CTSPP_72;
wire CTS_n333;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_21), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_21), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_21), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_21), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_21), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_21), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_21), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_21), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_21), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_21), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_21), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_21), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_21), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_21), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n333), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n333), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n333), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n333), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n333), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n333), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n333), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n333), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n333), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n333), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n333), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n333), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n333), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n333), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n333), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n333), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n333), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n333), .D (in[31]));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n333), .D (in[32]));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n333), .D (in[33]));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n333), .D (in[34]));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n333), .D (in[35]));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n333), .D (in[36]));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n333), .D (in[37]));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n333), .D (in[38]));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n333), .D (in[39]));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n333), .D (in[40]));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (clk_CTSPP_62), .D (in[41]));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (clk_CTSPP_62), .D (in[42]));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (clk_CTSPP_62), .D (in[43]));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (clk_CTSPP_62), .D (in[44]));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (clk_CTSPP_62), .D (in[45]));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (clk_CTSPP_62), .D (in[46]));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (clk_CTSPP_62), .D (in[47]));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (clk_CTSPP_62), .D (in[48]));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (clk_CTSPP_62), .D (in[49]));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (clk_CTSPP_62), .D (in[50]));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (clk_CTSPP_62), .D (in[51]));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (clk_CTSPP_62), .D (in[52]));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (clk_CTSPP_62), .D (in[53]));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (clk_CTSPP_62), .D (in[54]));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (clk_CTSPP_62), .D (in[55]));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (clk_CTSPP_62), .D (in[56]));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (clk_CTSPP_62), .D (in[57]));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (clk_CTSPP_62), .D (in[58]));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (clk_CTSPP_62), .D (in[59]));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (clk_CTSPP_62), .D (in[60]));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (clk_CTSPP_62), .D (in[61]));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (clk_CTSPP_62), .D (in[62]));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (clk_CTSPP_62), .D (in[63]));
CLKBUF_X2 CTS_L2_c15 (.Z (CTS_n333), .A (clk_CTSPP_72));

endmodule //Register__parameterized0

module Register (clk_CTSPP_48, clk_CTSPP_61, clk_CTSPP_70, in, clk, out);

output [31:0] out;
output clk_CTSPP_48;
output clk_CTSPP_61;
input clk;
input [31:0] in;
input clk_CTSPP_70;
wire drc_ipo_n6;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_48), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_48), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_48), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_48), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_48), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_48), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_48), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_48), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_48), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_48), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_48), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_48), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_48), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_48), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk_CTSPP_48), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk_CTSPP_48), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk_CTSPP_48), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk_CTSPP_48), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk_CTSPP_48), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk_CTSPP_48), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk_CTSPP_48), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk_CTSPP_48), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk_CTSPP_61), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk_CTSPP_61), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk_CTSPP_61), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk_CTSPP_61), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk_CTSPP_61), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk_CTSPP_61), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk_CTSPP_61), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk_CTSPP_61), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk_CTSPP_61), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (clk_CTSPP_48), .D (in[31]));
BUF_X4 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X2 CTS_L2_c28 (.Z (clk_CTSPP_61), .A (clk_CTSPP_70));
CLKBUF_X3 CTS_L2_c14 (.Z (clk_CTSPP_48), .A (clk_CTSPP_70));

endmodule //Register

module Register__5_0 (clk_CTSPP_23, clk_CTSPP_52, clk_CTSPP_60, in, clk, out);

output [31:0] out;
output clk_CTSPP_23;
input clk;
input [31:0] in;
input clk_CTSPP_52;
input clk_CTSPP_60;
wire drc_ipo_n6;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk_CTSPP_23), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk_CTSPP_23), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk_CTSPP_23), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk_CTSPP_23), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk_CTSPP_23), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk_CTSPP_23), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk_CTSPP_52), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk_CTSPP_23), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk_CTSPP_23), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk_CTSPP_23), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk_CTSPP_23), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk_CTSPP_23), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk_CTSPP_52), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk_CTSPP_23), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk_CTSPP_23), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk_CTSPP_23), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk_CTSPP_52), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk_CTSPP_23), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk_CTSPP_52), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk_CTSPP_52), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk_CTSPP_52), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk_CTSPP_23), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk_CTSPP_23), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk_CTSPP_23), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk_CTSPP_52), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk_CTSPP_52), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk_CTSPP_52), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk_CTSPP_52), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk_CTSPP_52), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk_CTSPP_52), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk_CTSPP_52), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (clk_CTSPP_52), .D (in[31]));
BUF_X8 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X3 CTS_L2_c9 (.Z (clk_CTSPP_23), .A (clk_CTSPP_60));

endmodule //Register__5_0

module datapath__0_38 (p_0, sum1);

output [63:0] p_0;
input [63:0] sum1;
wire n_0;
wire n_1;
wire n_173;
wire n_2;
wire n_175;
wire n_3;
wire n_171;
wire n_4;
wire n_5;
wire n_169;
wire n_6;
wire n_7;
wire n_167;
wire n_8;
wire n_9;
wire n_165;
wire n_10;
wire n_11;
wire n_163;
wire n_12;
wire n_13;
wire n_161;
wire n_14;
wire n_15;
wire n_159;
wire n_16;
wire n_17;
wire n_157;
wire n_18;
wire n_19;
wire n_155;
wire n_20;
wire n_21;
wire n_153;
wire n_22;
wire n_23;
wire n_151;
wire n_24;
wire n_25;
wire n_149;
wire n_26;
wire n_27;
wire n_147;
wire n_28;
wire n_29;
wire n_145;
wire n_30;
wire n_31;
wire n_143;
wire n_32;
wire n_33;
wire n_141;
wire n_34;
wire n_35;
wire n_139;
wire n_36;
wire n_37;
wire n_137;
wire n_38;
wire n_39;
wire n_135;
wire n_40;
wire n_41;
wire n_224;
wire n_42;
wire n_43;
wire n_223;
wire n_44;
wire n_45;
wire n_221;
wire n_46;
wire n_47;
wire n_219;
wire n_48;
wire n_49;
wire n_218;
wire n_50;
wire n_51;
wire n_216;
wire n_52;
wire n_53;
wire n_215;
wire n_54;
wire n_55;
wire n_214;
wire n_56;
wire n_57;
wire n_58;
wire n_213;
wire n_225;
wire n_59;
wire n_212;
wire n_60;
wire n_211;
wire n_226;
wire n_61;
wire n_209;
wire n_62;
wire n_210;
wire n_63;
wire n_190;
wire n_64;
wire n_65;
wire n_208;
wire n_66;
wire n_67;
wire n_71;
wire n_68;
wire n_69;
wire n_74;
wire n_189;
wire n_70;
wire n_207;
wire n_228;
wire n_72;
wire n_73;
wire n_206;
wire n_75;
wire n_76;
wire n_205;
wire n_229;
wire n_77;
wire n_204;
wire n_78;
wire n_187;
wire n_231;
wire n_79;
wire n_80;
wire n_202;
wire n_81;
wire n_185;
wire n_184;
wire n_82;
wire n_84;
wire n_233;
wire n_83;
wire n_199;
wire n_183;
wire n_86;
wire n_92;
wire n_87;
wire n_200;
wire n_88;
wire n_89;
wire n_90;
wire n_133;
wire n_91;
wire n_132;
wire n_131;
wire n_130;
wire n_93;
wire n_97;
wire n_94;
wire n_102;
wire n_95;
wire n_96;
wire n_100;
wire n_101;
wire n_127;
wire n_98;
wire n_181;
wire n_99;
wire n_128;
wire n_234;
wire n_103;
wire n_107;
wire n_104;
wire n_182;
wire n_105;
wire n_110;
wire n_106;
wire n_237;
wire n_236;
wire n_108;
wire n_109;
wire n_180;
wire n_124;
wire n_111;
wire n_123;
wire n_112;
wire n_113;
wire n_118;
wire n_122;
wire n_179;
wire n_114;
wire n_115;
wire n_121;
wire n_195;
wire n_116;
wire n_120;
wire n_117;
wire n_119;
wire n_177;
wire n_176;
wire n_178;
wire n_238;
wire n_126;
wire n_125;
wire n_129;
wire n_134;
wire n_136;
wire n_138;
wire n_140;
wire n_142;
wire n_144;
wire n_146;
wire n_148;
wire n_150;
wire n_152;
wire n_154;
wire n_156;
wire n_158;
wire n_160;
wire n_162;
wire n_164;
wire n_166;
wire n_168;
wire n_170;
wire n_172;
wire n_174;
wire n_197;
wire n_235;
wire n_186;
wire n_188;
wire n_203;
wire n_230;
wire n_191;
wire n_193;
wire n_192;
wire n_196;
wire n_198;
wire n_232;
wire n_201;
wire n_227;
wire n_217;
wire n_220;
wire n_222;


INV_X1 i_301 (.ZN (n_238), .A (sum1[58]));
INV_X1 i_300 (.ZN (n_237), .A (sum1[57]));
INV_X1 i_299 (.ZN (n_236), .A (sum1[56]));
INV_X1 i_298 (.ZN (n_235), .A (n_125));
INV_X1 i_297 (.ZN (n_234), .A (n_129));
INV_X1 i_296 (.ZN (n_233), .A (sum1[46]));
NOR3_X1 i_295 (.ZN (n_232), .A1 (sum1[45]), .A2 (sum1[47]), .A3 (sum1[44]));
INV_X1 i_294 (.ZN (n_231), .A (sum1[43]));
INV_X1 i_293 (.ZN (n_230), .A (sum1[42]));
INV_X1 i_292 (.ZN (n_229), .A (sum1[41]));
INV_X1 i_291 (.ZN (n_228), .A (sum1[37]));
NOR2_X1 i_290 (.ZN (n_227), .A1 (sum1[39]), .A2 (sum1[38]));
INV_X1 i_289 (.ZN (n_226), .A (sum1[33]));
INV_X1 i_288 (.ZN (n_225), .A (sum1[31]));
INV_X1 i_287 (.ZN (n_224), .A (n_134));
OR2_X1 i_286 (.ZN (n_223), .A1 (sum1[23]), .A2 (n_224));
NOR2_X1 i_285 (.ZN (n_222), .A1 (n_223), .A2 (sum1[24]));
INV_X1 i_284 (.ZN (n_221), .A (n_222));
NOR2_X1 i_283 (.ZN (n_220), .A1 (sum1[25]), .A2 (n_221));
INV_X1 i_282 (.ZN (n_219), .A (n_220));
OR2_X1 i_281 (.ZN (n_218), .A1 (sum1[26]), .A2 (n_219));
NOR2_X1 i_280 (.ZN (n_217), .A1 (sum1[27]), .A2 (n_218));
INV_X1 i_279 (.ZN (n_216), .A (n_217));
OR2_X1 i_278 (.ZN (n_215), .A1 (n_216), .A2 (sum1[28]));
OR2_X1 i_277 (.ZN (n_214), .A1 (n_215), .A2 (sum1[29]));
NOR2_X1 i_276 (.ZN (n_213), .A1 (n_214), .A2 (sum1[30]));
NAND2_X1 i_275 (.ZN (n_212), .A1 (n_225), .A2 (n_213));
NOR2_X1 i_274 (.ZN (n_211), .A1 (sum1[32]), .A2 (n_212));
NAND2_X1 i_273 (.ZN (n_210), .A1 (n_211), .A2 (n_226));
OR2_X1 i_272 (.ZN (n_209), .A1 (sum1[34]), .A2 (n_210));
OR3_X1 i_271 (.ZN (n_208), .A1 (n_209), .A2 (sum1[35]), .A3 (sum1[36]));
INV_X1 i_270 (.ZN (n_207), .A (n_208));
NAND3_X1 i_269 (.ZN (n_206), .A1 (n_207), .A2 (n_228), .A3 (n_227));
NOR2_X1 i_268 (.ZN (n_205), .A1 (n_206), .A2 (sum1[40]));
NAND2_X1 i_267 (.ZN (n_204), .A1 (n_205), .A2 (n_229));
INV_X1 i_266 (.ZN (n_203), .A (n_204));
NAND3_X1 i_265 (.ZN (n_202), .A1 (n_203), .A2 (n_231), .A3 (n_230));
INV_X1 i_264 (.ZN (n_201), .A (n_202));
NAND3_X1 i_263 (.ZN (n_200), .A1 (n_233), .A2 (n_232), .A3 (n_201));
INV_X1 i_262 (.ZN (n_199), .A (n_200));
NAND4_X1 i_261 (.ZN (n_198), .A1 (n_235), .A2 (n_234), .A3 (n_236), .A4 (n_199));
INV_X1 i_260 (.ZN (n_197), .A (n_198));
NOR2_X1 i_259 (.ZN (n_196), .A1 (sum1[59]), .A2 (sum1[60]));
NAND4_X1 i_258 (.ZN (n_195), .A1 (n_196), .A2 (n_197), .A3 (n_238), .A4 (n_237));
NAND2_X1 i_256 (.ZN (n_193), .A1 (n_176), .A2 (n_118));
NAND2_X1 i_255 (.ZN (n_192), .A1 (sum1[61]), .A2 (n_195));
NAND2_X1 i_254 (.ZN (n_191), .A1 (n_193), .A2 (n_192));
INV_X1 i_253 (.ZN (p_0[61]), .A (n_191));
OR2_X1 i_252 (.ZN (n_190), .A1 (n_209), .A2 (sum1[35]));
INV_X1 i_251 (.ZN (n_189), .A (sum1[38]));
NAND2_X1 i_250 (.ZN (n_188), .A1 (n_203), .A2 (n_230));
INV_X1 i_249 (.ZN (n_187), .A (n_188));
OR2_X1 i_248 (.ZN (n_186), .A1 (n_202), .A2 (sum1[44]));
INV_X1 i_247 (.ZN (n_185), .A (n_186));
INV_X1 i_246 (.ZN (n_184), .A (sum1[45]));
INV_X1 i_245 (.ZN (n_183), .A (sum1[47]));
NAND3_X2 i_244 (.ZN (n_182), .A1 (n_235), .A2 (n_234), .A3 (n_199));
INV_X2 i_243 (.ZN (n_181), .A (n_182));
NAND3_X1 i_242 (.ZN (n_180), .A1 (n_197), .A2 (n_238), .A3 (n_237));
INV_X1 i_241 (.ZN (n_179), .A (sum1[60]));
INV_X1 i_240 (.ZN (n_178), .A (sum1[59]));
INV_X1 i_239 (.ZN (n_177), .A (sum1[62]));
INV_X1 i_238 (.ZN (n_176), .A (sum1[61]));
OR2_X1 i_237 (.ZN (n_175), .A1 (sum1[1]), .A2 (sum1[0]));
NOR2_X1 i_236 (.ZN (n_174), .A1 (sum1[2]), .A2 (n_175));
INV_X1 i_235 (.ZN (n_173), .A (n_174));
NOR2_X1 i_234 (.ZN (n_172), .A1 (sum1[3]), .A2 (n_173));
INV_X1 i_233 (.ZN (n_171), .A (n_172));
NOR2_X1 i_232 (.ZN (n_170), .A1 (sum1[4]), .A2 (n_171));
INV_X1 i_231 (.ZN (n_169), .A (n_170));
NOR2_X1 i_230 (.ZN (n_168), .A1 (sum1[5]), .A2 (n_169));
INV_X1 i_229 (.ZN (n_167), .A (n_168));
NOR2_X1 i_228 (.ZN (n_166), .A1 (sum1[6]), .A2 (n_167));
INV_X1 i_227 (.ZN (n_165), .A (n_166));
NOR2_X1 i_226 (.ZN (n_164), .A1 (sum1[7]), .A2 (n_165));
INV_X1 i_225 (.ZN (n_163), .A (n_164));
NOR2_X1 i_224 (.ZN (n_162), .A1 (sum1[8]), .A2 (n_163));
INV_X1 i_223 (.ZN (n_161), .A (n_162));
NOR2_X1 i_222 (.ZN (n_160), .A1 (sum1[9]), .A2 (n_161));
INV_X1 i_221 (.ZN (n_159), .A (n_160));
NOR2_X1 i_220 (.ZN (n_158), .A1 (sum1[10]), .A2 (n_159));
INV_X1 i_219 (.ZN (n_157), .A (n_158));
NOR2_X1 i_218 (.ZN (n_156), .A1 (sum1[11]), .A2 (n_157));
INV_X1 i_217 (.ZN (n_155), .A (n_156));
NOR2_X1 i_216 (.ZN (n_154), .A1 (sum1[12]), .A2 (n_155));
INV_X1 i_215 (.ZN (n_153), .A (n_154));
NOR2_X1 i_214 (.ZN (n_152), .A1 (sum1[13]), .A2 (n_153));
INV_X1 i_213 (.ZN (n_151), .A (n_152));
NOR2_X1 i_212 (.ZN (n_150), .A1 (sum1[14]), .A2 (n_151));
INV_X1 i_211 (.ZN (n_149), .A (n_150));
NOR2_X1 i_210 (.ZN (n_148), .A1 (sum1[15]), .A2 (n_149));
INV_X1 i_209 (.ZN (n_147), .A (n_148));
NOR2_X1 i_208 (.ZN (n_146), .A1 (sum1[16]), .A2 (n_147));
INV_X1 i_207 (.ZN (n_145), .A (n_146));
NOR2_X1 i_206 (.ZN (n_144), .A1 (sum1[17]), .A2 (n_145));
INV_X1 i_205 (.ZN (n_143), .A (n_144));
NOR2_X1 i_204 (.ZN (n_142), .A1 (sum1[18]), .A2 (n_143));
INV_X1 i_203 (.ZN (n_141), .A (n_142));
NOR2_X1 i_202 (.ZN (n_140), .A1 (sum1[19]), .A2 (n_141));
INV_X1 i_201 (.ZN (n_139), .A (n_140));
NOR2_X1 i_200 (.ZN (n_138), .A1 (sum1[20]), .A2 (n_139));
INV_X1 i_199 (.ZN (n_137), .A (n_138));
NOR2_X1 i_198 (.ZN (n_136), .A1 (sum1[21]), .A2 (n_137));
INV_X1 i_197 (.ZN (n_135), .A (n_136));
NOR2_X1 i_196 (.ZN (n_134), .A1 (sum1[22]), .A2 (n_135));
INV_X1 i_195 (.ZN (n_133), .A (sum1[51]));
INV_X1 i_194 (.ZN (n_132), .A (sum1[50]));
INV_X1 i_193 (.ZN (n_131), .A (sum1[49]));
INV_X1 i_192 (.ZN (n_130), .A (sum1[48]));
NAND4_X1 i_191 (.ZN (n_129), .A1 (n_132), .A2 (n_131), .A3 (n_133), .A4 (n_130));
INV_X1 i_190 (.ZN (n_128), .A (sum1[53]));
INV_X1 i_189 (.ZN (n_127), .A (sum1[52]));
NOR2_X2 i_188 (.ZN (n_126), .A1 (sum1[54]), .A2 (sum1[55]));
NAND3_X1 i_187 (.ZN (n_125), .A1 (n_128), .A2 (n_127), .A3 (n_126));
NOR2_X1 i_186 (.ZN (n_124), .A1 (sum1[57]), .A2 (sum1[56]));
NAND4_X1 i_185 (.ZN (n_123), .A1 (n_124), .A2 (n_178), .A3 (n_238), .A4 (n_181));
INV_X1 i_184 (.ZN (n_122), .A (n_123));
NAND4_X1 i_183 (.ZN (n_121), .A1 (n_122), .A2 (n_177), .A3 (n_176), .A4 (n_179));
NAND2_X1 i_182 (.ZN (n_120), .A1 (n_121), .A2 (sum1[63]));
INV_X1 i_181 (.ZN (n_119), .A (sum1[63]));
INV_X1 i_180 (.ZN (n_118), .A (n_195));
NAND4_X1 i_179 (.ZN (n_117), .A1 (n_118), .A2 (n_119), .A3 (n_177), .A4 (n_176));
NAND2_X1 i_178 (.ZN (n_116), .A1 (n_120), .A2 (n_117));
INV_X1 i_177 (.ZN (p_0[63]), .A (n_116));
OAI21_X1 i_176 (.ZN (n_115), .A (sum1[62]), .B1 (n_195), .B2 (sum1[61]));
NAND2_X1 i_175 (.ZN (n_114), .A1 (n_115), .A2 (n_121));
INV_X1 i_174 (.ZN (p_0[62]), .A (n_114));
NOR2_X1 i_173 (.ZN (n_113), .A1 (n_122), .A2 (n_179));
NOR2_X1 i_172 (.ZN (p_0[60]), .A1 (n_113), .A2 (n_118));
NAND2_X1 i_171 (.ZN (n_112), .A1 (n_180), .A2 (sum1[59]));
NAND2_X1 i_170 (.ZN (n_111), .A1 (n_123), .A2 (n_112));
INV_X1 i_169 (.ZN (p_0[59]), .A (n_111));
NAND2_X1 i_168 (.ZN (n_110), .A1 (n_124), .A2 (n_181));
NAND2_X1 i_167 (.ZN (n_109), .A1 (n_110), .A2 (sum1[58]));
NAND2_X1 i_166 (.ZN (n_108), .A1 (n_109), .A2 (n_180));
INV_X1 i_165 (.ZN (p_0[58]), .A (n_108));
NAND2_X1 i_164 (.ZN (n_107), .A1 (n_181), .A2 (n_236));
INV_X1 i_163 (.ZN (n_106), .A (n_107));
OAI21_X1 i_162 (.ZN (n_105), .A (n_110), .B1 (n_106), .B2 (n_237));
INV_X1 i_161 (.ZN (p_0[57]), .A (n_105));
NAND2_X1 i_160 (.ZN (n_104), .A1 (n_182), .A2 (sum1[56]));
NAND2_X1 i_159 (.ZN (n_103), .A1 (n_107), .A2 (n_104));
INV_X1 i_158 (.ZN (p_0[56]), .A (n_103));
NAND2_X1 i_157 (.ZN (n_102), .A1 (n_199), .A2 (n_234));
INV_X1 i_156 (.ZN (n_101), .A (n_102));
NAND3_X1 i_155 (.ZN (n_100), .A1 (n_101), .A2 (n_128), .A3 (n_127));
OR2_X1 i_154 (.ZN (n_99), .A1 (n_100), .A2 (sum1[54]));
AOI21_X1 i_153 (.ZN (p_0[55]), .A (n_181), .B1 (n_99), .B2 (sum1[55]));
XNOR2_X1 i_152 (.ZN (n_98), .A (n_100), .B (sum1[54]));
INV_X1 i_151 (.ZN (p_0[54]), .A (n_98));
NAND2_X1 i_150 (.ZN (n_97), .A1 (n_101), .A2 (n_127));
NAND2_X1 i_149 (.ZN (n_96), .A1 (n_97), .A2 (sum1[53]));
NAND2_X1 i_148 (.ZN (n_95), .A1 (n_96), .A2 (n_100));
INV_X1 i_147 (.ZN (p_0[53]), .A (n_95));
NAND2_X1 i_146 (.ZN (n_94), .A1 (n_102), .A2 (sum1[52]));
NAND2_X1 i_145 (.ZN (n_93), .A1 (n_97), .A2 (n_94));
INV_X1 i_144 (.ZN (p_0[52]), .A (n_93));
NAND2_X1 i_143 (.ZN (n_92), .A1 (n_199), .A2 (n_130));
INV_X1 i_142 (.ZN (n_91), .A (n_92));
NAND3_X1 i_141 (.ZN (n_90), .A1 (n_91), .A2 (n_132), .A3 (n_131));
XNOR2_X1 i_140 (.ZN (p_0[51]), .A (n_90), .B (n_133));
OAI21_X1 i_139 (.ZN (n_89), .A (sum1[50]), .B1 (n_92), .B2 (sum1[49]));
AND2_X1 i_138 (.ZN (p_0[50]), .A1 (n_89), .A2 (n_90));
XNOR2_X1 i_137 (.ZN (n_88), .A (n_92), .B (sum1[49]));
INV_X1 i_136 (.ZN (p_0[49]), .A (n_88));
NAND2_X1 i_135 (.ZN (n_87), .A1 (n_200), .A2 (sum1[48]));
NAND2_X1 i_134 (.ZN (n_86), .A1 (n_92), .A2 (n_87));
INV_X1 i_133 (.ZN (p_0[48]), .A (n_86));
NOR2_X1 i_131 (.ZN (n_84), .A1 (n_186), .A2 (sum1[45]));
AOI21_X1 i_130 (.ZN (n_83), .A (n_183), .B1 (n_84), .B2 (n_233));
NOR2_X1 i_129 (.ZN (p_0[47]), .A1 (n_83), .A2 (n_199));
XNOR2_X1 i_128 (.ZN (n_82), .A (n_84), .B (n_233));
INV_X1 i_127 (.ZN (p_0[46]), .A (n_82));
XNOR2_X1 i_126 (.ZN (n_81), .A (n_185), .B (n_184));
INV_X1 i_125 (.ZN (p_0[45]), .A (n_81));
NAND2_X1 i_124 (.ZN (n_80), .A1 (n_202), .A2 (sum1[44]));
NAND2_X1 i_123 (.ZN (n_79), .A1 (n_186), .A2 (n_80));
INV_X1 i_122 (.ZN (p_0[44]), .A (n_79));
XNOR2_X1 i_121 (.ZN (n_78), .A (n_187), .B (n_231));
INV_X1 i_120 (.ZN (p_0[43]), .A (n_78));
XNOR2_X1 i_119 (.ZN (n_77), .A (n_204), .B (sum1[42]));
INV_X1 i_118 (.ZN (p_0[42]), .A (n_77));
XNOR2_X1 i_117 (.ZN (n_76), .A (n_205), .B (n_229));
INV_X1 i_116 (.ZN (p_0[41]), .A (n_76));
XNOR2_X1 i_115 (.ZN (n_75), .A (sum1[40]), .B (n_206));
INV_X1 i_114 (.ZN (p_0[40]), .A (n_75));
NAND3_X1 i_113 (.ZN (n_74), .A1 (n_207), .A2 (n_189), .A3 (n_228));
NAND2_X1 i_112 (.ZN (n_73), .A1 (n_74), .A2 (sum1[39]));
NAND2_X1 i_111 (.ZN (n_72), .A1 (n_73), .A2 (n_206));
INV_X1 i_110 (.ZN (p_0[39]), .A (n_72));
NAND2_X1 i_109 (.ZN (n_71), .A1 (n_207), .A2 (n_228));
INV_X1 i_108 (.ZN (n_70), .A (n_71));
OAI21_X1 i_107 (.ZN (n_69), .A (n_74), .B1 (n_189), .B2 (n_70));
INV_X1 i_106 (.ZN (p_0[38]), .A (n_69));
NAND2_X1 i_105 (.ZN (n_68), .A1 (n_208), .A2 (sum1[37]));
NAND2_X1 i_104 (.ZN (n_67), .A1 (n_71), .A2 (n_68));
INV_X1 i_103 (.ZN (p_0[37]), .A (n_67));
NAND2_X1 i_102 (.ZN (n_66), .A1 (n_190), .A2 (sum1[36]));
NAND2_X1 i_101 (.ZN (n_65), .A1 (n_208), .A2 (n_66));
INV_X1 i_100 (.ZN (p_0[36]), .A (n_65));
NAND2_X1 i_99 (.ZN (n_64), .A1 (n_209), .A2 (sum1[35]));
NAND2_X1 i_98 (.ZN (n_63), .A1 (n_190), .A2 (n_64));
INV_X1 i_97 (.ZN (p_0[35]), .A (n_63));
NAND2_X1 i_96 (.ZN (n_62), .A1 (n_210), .A2 (sum1[34]));
NAND2_X1 i_95 (.ZN (n_61), .A1 (n_209), .A2 (n_62));
INV_X1 i_94 (.ZN (p_0[34]), .A (n_61));
XNOR2_X1 i_93 (.ZN (n_60), .A (n_211), .B (n_226));
INV_X1 i_92 (.ZN (p_0[33]), .A (n_60));
XNOR2_X1 i_91 (.ZN (n_59), .A (sum1[32]), .B (n_212));
INV_X1 i_90 (.ZN (p_0[32]), .A (n_59));
XNOR2_X1 i_89 (.ZN (n_58), .A (n_213), .B (n_225));
INV_X1 i_88 (.ZN (p_0[31]), .A (n_58));
XNOR2_X1 i_87 (.ZN (n_57), .A (sum1[30]), .B (n_214));
INV_X1 i_86 (.ZN (p_0[30]), .A (n_57));
NAND2_X1 i_85 (.ZN (n_56), .A1 (sum1[29]), .A2 (n_215));
NAND2_X1 i_84 (.ZN (n_55), .A1 (n_214), .A2 (n_56));
INV_X1 i_83 (.ZN (p_0[29]), .A (n_55));
NAND2_X1 i_82 (.ZN (n_54), .A1 (n_216), .A2 (sum1[28]));
NAND2_X1 i_81 (.ZN (n_53), .A1 (n_215), .A2 (n_54));
INV_X1 i_80 (.ZN (p_0[28]), .A (n_53));
NAND2_X1 i_79 (.ZN (n_52), .A1 (sum1[27]), .A2 (n_218));
NAND2_X1 i_78 (.ZN (n_51), .A1 (n_216), .A2 (n_52));
INV_X1 i_77 (.ZN (p_0[27]), .A (n_51));
NAND2_X1 i_76 (.ZN (n_50), .A1 (sum1[26]), .A2 (n_219));
NAND2_X1 i_75 (.ZN (n_49), .A1 (n_218), .A2 (n_50));
INV_X1 i_74 (.ZN (p_0[26]), .A (n_49));
NAND2_X1 i_73 (.ZN (n_48), .A1 (sum1[25]), .A2 (n_221));
NAND2_X1 i_72 (.ZN (n_47), .A1 (n_219), .A2 (n_48));
INV_X1 i_71 (.ZN (p_0[25]), .A (n_47));
NAND2_X1 i_70 (.ZN (n_46), .A1 (sum1[24]), .A2 (n_223));
NAND2_X1 i_69 (.ZN (n_45), .A1 (n_221), .A2 (n_46));
INV_X1 i_68 (.ZN (p_0[24]), .A (n_45));
NAND2_X1 i_67 (.ZN (n_44), .A1 (sum1[23]), .A2 (n_224));
NAND2_X1 i_66 (.ZN (n_43), .A1 (n_223), .A2 (n_44));
INV_X1 i_65 (.ZN (p_0[23]), .A (n_43));
NAND2_X1 i_64 (.ZN (n_42), .A1 (sum1[22]), .A2 (n_135));
NAND2_X1 i_63 (.ZN (n_41), .A1 (n_224), .A2 (n_42));
INV_X1 i_62 (.ZN (p_0[22]), .A (n_41));
NAND2_X1 i_61 (.ZN (n_40), .A1 (sum1[21]), .A2 (n_137));
NAND2_X1 i_60 (.ZN (n_39), .A1 (n_135), .A2 (n_40));
INV_X1 i_59 (.ZN (p_0[21]), .A (n_39));
NAND2_X1 i_58 (.ZN (n_38), .A1 (sum1[20]), .A2 (n_139));
NAND2_X1 i_57 (.ZN (n_37), .A1 (n_137), .A2 (n_38));
INV_X1 i_56 (.ZN (p_0[20]), .A (n_37));
NAND2_X1 i_55 (.ZN (n_36), .A1 (sum1[19]), .A2 (n_141));
NAND2_X1 i_54 (.ZN (n_35), .A1 (n_139), .A2 (n_36));
INV_X1 i_53 (.ZN (p_0[19]), .A (n_35));
NAND2_X1 i_52 (.ZN (n_34), .A1 (sum1[18]), .A2 (n_143));
NAND2_X1 i_51 (.ZN (n_33), .A1 (n_141), .A2 (n_34));
INV_X1 i_50 (.ZN (p_0[18]), .A (n_33));
NAND2_X1 i_49 (.ZN (n_32), .A1 (sum1[17]), .A2 (n_145));
NAND2_X1 i_48 (.ZN (n_31), .A1 (n_143), .A2 (n_32));
INV_X1 i_47 (.ZN (p_0[17]), .A (n_31));
NAND2_X1 i_46 (.ZN (n_30), .A1 (sum1[16]), .A2 (n_147));
NAND2_X1 i_45 (.ZN (n_29), .A1 (n_145), .A2 (n_30));
INV_X1 i_44 (.ZN (p_0[16]), .A (n_29));
NAND2_X1 i_43 (.ZN (n_28), .A1 (sum1[15]), .A2 (n_149));
NAND2_X1 i_42 (.ZN (n_27), .A1 (n_147), .A2 (n_28));
INV_X1 i_41 (.ZN (p_0[15]), .A (n_27));
NAND2_X1 i_40 (.ZN (n_26), .A1 (sum1[14]), .A2 (n_151));
NAND2_X1 i_39 (.ZN (n_25), .A1 (n_149), .A2 (n_26));
INV_X1 i_38 (.ZN (p_0[14]), .A (n_25));
NAND2_X1 i_37 (.ZN (n_24), .A1 (sum1[13]), .A2 (n_153));
NAND2_X1 i_36 (.ZN (n_23), .A1 (n_151), .A2 (n_24));
INV_X1 i_35 (.ZN (p_0[13]), .A (n_23));
NAND2_X1 i_34 (.ZN (n_22), .A1 (sum1[12]), .A2 (n_155));
NAND2_X1 i_33 (.ZN (n_21), .A1 (n_153), .A2 (n_22));
INV_X1 i_32 (.ZN (p_0[12]), .A (n_21));
NAND2_X1 i_31 (.ZN (n_20), .A1 (sum1[11]), .A2 (n_157));
NAND2_X1 i_30 (.ZN (n_19), .A1 (n_155), .A2 (n_20));
INV_X1 i_29 (.ZN (p_0[11]), .A (n_19));
NAND2_X1 i_28 (.ZN (n_18), .A1 (sum1[10]), .A2 (n_159));
NAND2_X1 i_27 (.ZN (n_17), .A1 (n_157), .A2 (n_18));
INV_X1 i_26 (.ZN (p_0[10]), .A (n_17));
NAND2_X1 i_25 (.ZN (n_16), .A1 (sum1[9]), .A2 (n_161));
NAND2_X1 i_24 (.ZN (n_15), .A1 (n_159), .A2 (n_16));
INV_X1 i_23 (.ZN (p_0[9]), .A (n_15));
NAND2_X1 i_22 (.ZN (n_14), .A1 (sum1[8]), .A2 (n_163));
NAND2_X1 i_21 (.ZN (n_13), .A1 (n_161), .A2 (n_14));
INV_X1 i_20 (.ZN (p_0[8]), .A (n_13));
NAND2_X1 i_19 (.ZN (n_12), .A1 (sum1[7]), .A2 (n_165));
NAND2_X1 i_18 (.ZN (n_11), .A1 (n_163), .A2 (n_12));
INV_X1 i_17 (.ZN (p_0[7]), .A (n_11));
NAND2_X1 i_16 (.ZN (n_10), .A1 (sum1[6]), .A2 (n_167));
NAND2_X1 i_15 (.ZN (n_9), .A1 (n_165), .A2 (n_10));
INV_X1 i_14 (.ZN (p_0[6]), .A (n_9));
NAND2_X1 i_13 (.ZN (n_8), .A1 (sum1[5]), .A2 (n_169));
NAND2_X1 i_12 (.ZN (n_7), .A1 (n_167), .A2 (n_8));
INV_X1 i_11 (.ZN (p_0[5]), .A (n_7));
NAND2_X1 i_10 (.ZN (n_6), .A1 (sum1[4]), .A2 (n_171));
NAND2_X1 i_9 (.ZN (n_5), .A1 (n_169), .A2 (n_6));
INV_X1 i_8 (.ZN (p_0[4]), .A (n_5));
NAND2_X1 i_7 (.ZN (n_4), .A1 (sum1[3]), .A2 (n_173));
NAND2_X1 i_6 (.ZN (n_3), .A1 (n_171), .A2 (n_4));
INV_X1 i_5 (.ZN (p_0[3]), .A (n_3));
NAND2_X1 i_4 (.ZN (n_2), .A1 (sum1[2]), .A2 (n_175));
NAND2_X1 i_3 (.ZN (n_1), .A1 (n_173), .A2 (n_2));
INV_X1 i_2 (.ZN (p_0[2]), .A (n_1));
XNOR2_X1 i_1 (.ZN (n_0), .A (sum1[1]), .B (sum1[0]));
INV_X1 i_0 (.ZN (p_0[1]), .A (n_0));

endmodule //datapath__0_38

module datapath__0_3 (p_0, a);

output [31:0] p_0;
input [31:0] a;
wire n_0;
wire n_4;
wire n_1;
wire n_2;
wire n_3;
wire n_7;
wire n_142;
wire n_143;
wire n_5;
wire n_6;
wire n_141;
wire n_144;
wire n_8;
wire n_13;
wire n_9;
wire n_10;
wire n_15;
wire n_104;
wire n_11;
wire n_12;
wire n_14;
wire n_125;
wire n_124;
wire n_16;
wire n_20;
wire n_17;
wire n_40;
wire n_18;
wire n_19;
wire n_21;
wire n_39;
wire n_128;
wire n_37;
wire n_129;
wire n_22;
wire n_31;
wire n_23;
wire n_38;
wire n_24;
wire n_25;
wire n_28;
wire n_26;
wire n_135;
wire n_27;
wire n_42;
wire n_134;
wire n_133;
wire n_29;
wire n_35;
wire n_138;
wire n_30;
wire n_41;
wire n_32;
wire n_33;
wire n_139;
wire n_34;
wire n_137;
wire n_36;
wire n_126;
wire n_140;
wire n_120;
wire n_43;
wire n_87;
wire n_44;
wire n_45;
wire n_46;
wire n_84;
wire n_86;
wire n_122;
wire n_108;
wire n_47;
wire n_48;
wire n_88;
wire n_85;
wire n_49;
wire n_51;
wire n_67;
wire n_81;
wire n_50;
wire n_55;
wire n_82;
wire n_52;
wire n_100;
wire n_53;
wire n_54;
wire n_56;
wire n_57;
wire n_63;
wire n_58;
wire n_80;
wire n_59;
wire n_60;
wire n_61;
wire n_64;
wire n_73;
wire n_75;
wire n_78;
wire n_62;
wire n_71;
wire n_65;
wire n_66;
wire n_69;
wire n_68;
wire n_99;
wire n_70;
wire n_72;
wire n_77;
wire n_74;
wire n_76;
wire n_79;
wire n_83;
wire n_146;
wire n_118;
wire n_89;
wire n_115;
wire n_90;
wire n_91;
wire n_95;
wire n_92;
wire n_97;
wire n_93;
wire n_94;
wire n_96;
wire n_116;
wire n_112;
wire n_105;
wire n_111;
wire n_101;
wire n_113;
wire n_107;
wire n_106;
wire n_109;
wire n_102;
wire n_110;
wire n_132;
wire n_114;
wire n_117;
wire n_119;
wire n_131;
wire n_121;
wire n_103;
wire n_127;
wire n_130;
wire n_145;
wire n_147;
wire n_123;


INV_X1 i_176 (.ZN (n_123), .A (a[18]));
INV_X1 i_175 (.ZN (n_122), .A (a[17]));
INV_X1 i_174 (.ZN (n_108), .A (a[16]));
NOR4_X1 i_172 (.ZN (n_107), .A1 (a[18]), .A2 (a[16]), .A3 (a[17]), .A4 (a[23]));
INV_X2 i_171 (.ZN (n_104), .A (a[5]));
INV_X1 i_170 (.ZN (n_103), .A (a[4]));
NOR2_X1 i_169 (.ZN (n_102), .A1 (a[5]), .A2 (a[4]));
NAND3_X1 i_178 (.ZN (n_147), .A1 (n_108), .A2 (n_123), .A3 (n_122));
INV_X1 i_177 (.ZN (n_146), .A (n_147));
INV_X1 i_168 (.ZN (n_145), .A (a[3]));
INV_X1 i_167 (.ZN (n_144), .A (a[2]));
INV_X1 i_166 (.ZN (n_143), .A (a[1]));
INV_X1 i_173 (.ZN (n_142), .A (a[0]));
NAND4_X2 i_165 (.ZN (n_141), .A1 (n_142), .A2 (n_145), .A3 (n_144), .A4 (n_143));
INV_X2 i_164 (.ZN (n_140), .A (n_141));
INV_X1 i_163 (.ZN (n_139), .A (a[15]));
INV_X1 i_162 (.ZN (n_138), .A (a[14]));
NAND2_X1 i_161 (.ZN (n_137), .A1 (n_139), .A2 (n_138));
INV_X1 i_159 (.ZN (n_135), .A (a[13]));
INV_X1 i_158 (.ZN (n_134), .A (a[12]));
INV_X2 i_157 (.ZN (n_133), .A (a[11]));
NAND3_X2 i_156 (.ZN (n_132), .A1 (n_134), .A2 (n_133), .A3 (n_135));
INV_X2 i_155 (.ZN (n_131), .A (n_132));
INV_X1 i_154 (.ZN (n_130), .A (a[10]));
INV_X2 i_153 (.ZN (n_129), .A (a[9]));
INV_X2 i_152 (.ZN (n_128), .A (a[8]));
NAND3_X1 i_151 (.ZN (n_127), .A1 (n_130), .A2 (n_129), .A3 (n_128));
INV_X2 i_150 (.ZN (n_126), .A (n_127));
INV_X2 i_149 (.ZN (n_125), .A (a[7]));
INV_X2 i_148 (.ZN (n_124), .A (a[6]));
NAND4_X2 i_147 (.ZN (n_121), .A1 (n_103), .A2 (n_104), .A3 (n_124), .A4 (n_125));
INV_X2 i_146 (.ZN (n_120), .A (n_121));
NAND4_X2 i_145 (.ZN (n_119), .A1 (n_120), .A2 (n_34), .A3 (n_131), .A4 (n_126));
INV_X4 i_144 (.ZN (n_118), .A (n_119));
INV_X1 i_141 (.ZN (n_117), .A (a[22]));
INV_X1 i_140 (.ZN (n_116), .A (a[20]));
INV_X1 i_139 (.ZN (n_115), .A (a[19]));
NAND4_X1 i_138 (.ZN (n_114), .A1 (n_83), .A2 (n_116), .A3 (n_115), .A4 (n_117));
INV_X1 i_137 (.ZN (n_113), .A (n_114));
NAND4_X1 i_143 (.ZN (n_112), .A1 (n_118), .A2 (n_146), .A3 (n_140), .A4 (n_113));
NOR2_X1 i_142 (.ZN (n_111), .A1 (n_132), .A2 (n_137));
NAND2_X1 i_136 (.ZN (n_110), .A1 (n_124), .A2 (n_125));
INV_X1 i_135 (.ZN (n_109), .A (n_110));
NAND3_X1 i_134 (.ZN (n_106), .A1 (n_126), .A2 (n_109), .A3 (n_102));
INV_X1 i_133 (.ZN (n_105), .A (n_106));
NAND2_X1 i_132 (.ZN (n_101), .A1 (n_113), .A2 (n_107));
INV_X2 i_131 (.ZN (n_100), .A (n_101));
NAND4_X1 i_130 (.ZN (n_99), .A1 (n_100), .A2 (n_105), .A3 (n_140), .A4 (n_111));
AOI21_X1 i_128 (.ZN (p_0[23]), .A (n_67), .B1 (n_112), .B2 (a[23]));
INV_X1 i_127 (.ZN (n_97), .A (n_112));
NAND2_X1 i_126 (.ZN (n_96), .A1 (n_116), .A2 (n_115));
INV_X1 i_125 (.ZN (n_95), .A (n_96));
NAND2_X1 i_124 (.ZN (n_94), .A1 (n_95), .A2 (n_83));
INV_X1 i_123 (.ZN (n_93), .A (n_94));
NAND4_X1 i_122 (.ZN (n_92), .A1 (n_118), .A2 (n_146), .A3 (n_140), .A4 (n_93));
AOI21_X1 i_121 (.ZN (p_0[22]), .A (n_97), .B1 (n_92), .B2 (a[22]));
INV_X1 i_120 (.ZN (n_91), .A (n_92));
NAND4_X1 i_119 (.ZN (n_90), .A1 (n_118), .A2 (n_146), .A3 (n_140), .A4 (n_95));
AOI21_X1 i_118 (.ZN (p_0[21]), .A (n_91), .B1 (n_90), .B2 (a[21]));
INV_X1 i_117 (.ZN (n_89), .A (n_90));
NAND4_X1 i_116 (.ZN (n_88), .A1 (n_118), .A2 (n_115), .A3 (n_146), .A4 (n_140));
AOI21_X1 i_115 (.ZN (p_0[20]), .A (n_89), .B1 (n_88), .B2 (a[20]));
NAND2_X2 i_114 (.ZN (n_87), .A1 (n_118), .A2 (n_140));
INV_X4 i_113 (.ZN (n_86), .A (n_87));
NAND2_X1 i_112 (.ZN (n_85), .A1 (n_86), .A2 (n_146));
INV_X1 i_111 (.ZN (n_84), .A (n_85));
INV_X1 i_110 (.ZN (n_83), .A (a[21]));
INV_X1 i_109 (.ZN (n_82), .A (a[25]));
INV_X1 i_108 (.ZN (n_81), .A (a[24]));
NAND2_X1 i_107 (.ZN (n_80), .A1 (n_82), .A2 (n_81));
OR3_X1 i_106 (.ZN (n_79), .A1 (n_80), .A2 (a[27]), .A3 (a[26]));
INV_X1 i_105 (.ZN (n_78), .A (n_79));
INV_X1 i_104 (.ZN (n_77), .A (a[30]));
INV_X1 i_103 (.ZN (n_76), .A (a[29]));
INV_X1 i_102 (.ZN (n_75), .A (a[28]));
NAND2_X1 i_101 (.ZN (n_74), .A1 (n_76), .A2 (n_75));
INV_X1 i_100 (.ZN (n_73), .A (n_74));
NAND2_X1 i_99 (.ZN (n_72), .A1 (n_73), .A2 (n_77));
INV_X1 i_98 (.ZN (n_71), .A (n_72));
NAND4_X1 i_97 (.ZN (n_70), .A1 (n_100), .A2 (n_86), .A3 (n_78), .A4 (n_71));
NAND2_X1 i_96 (.ZN (n_69), .A1 (n_70), .A2 (a[31]));
INV_X1 i_95 (.ZN (n_68), .A (a[31]));
INV_X2 i_94 (.ZN (n_67), .A (n_99));
NAND4_X1 i_93 (.ZN (n_66), .A1 (n_67), .A2 (n_68), .A3 (n_78), .A4 (n_71));
NAND2_X1 i_92 (.ZN (n_65), .A1 (n_66), .A2 (n_69));
INV_X1 i_91 (.ZN (p_0[31]), .A (n_65));
NAND3_X2 i_90 (.ZN (n_64), .A1 (n_100), .A2 (n_86), .A3 (n_78));
INV_X2 i_89 (.ZN (n_63), .A (n_64));
NAND4_X1 i_88 (.ZN (n_62), .A1 (n_100), .A2 (n_86), .A3 (n_78), .A4 (n_73));
AOI22_X1 i_87 (.ZN (p_0[30]), .A1 (n_62), .A2 (a[30]), .B1 (n_63), .B2 (n_71));
NAND4_X1 i_86 (.ZN (n_61), .A1 (n_100), .A2 (n_86), .A3 (n_75), .A4 (n_78));
AOI22_X1 i_85 (.ZN (p_0[29]), .A1 (n_61), .A2 (a[29]), .B1 (n_63), .B2 (n_73));
NAND2_X1 i_84 (.ZN (n_60), .A1 (n_64), .A2 (a[28]));
NAND2_X1 i_83 (.ZN (n_59), .A1 (n_60), .A2 (n_61));
INV_X1 i_82 (.ZN (p_0[28]), .A (n_59));
INV_X1 i_81 (.ZN (n_58), .A (a[26]));
INV_X1 i_80 (.ZN (n_57), .A (n_80));
NAND4_X1 i_79 (.ZN (n_56), .A1 (n_100), .A2 (n_86), .A3 (n_58), .A4 (n_57));
AOI21_X1 i_78 (.ZN (p_0[27]), .A (n_63), .B1 (n_56), .B2 (a[27]));
NAND3_X1 i_77 (.ZN (n_55), .A1 (n_100), .A2 (n_86), .A3 (n_57));
NAND2_X1 i_76 (.ZN (n_54), .A1 (n_55), .A2 (a[26]));
NAND2_X1 i_75 (.ZN (n_53), .A1 (n_54), .A2 (n_56));
INV_X1 i_74 (.ZN (p_0[26]), .A (n_53));
NAND3_X1 i_73 (.ZN (n_52), .A1 (n_100), .A2 (n_86), .A3 (n_81));
INV_X1 i_72 (.ZN (n_51), .A (n_52));
OAI21_X1 i_71 (.ZN (n_50), .A (n_55), .B1 (n_51), .B2 (n_82));
INV_X1 i_70 (.ZN (p_0[25]), .A (n_50));
NOR2_X1 i_69 (.ZN (n_49), .A1 (n_67), .A2 (n_81));
NOR2_X1 i_68 (.ZN (p_0[24]), .A1 (n_49), .A2 (n_51));
NAND2_X1 i_67 (.ZN (n_48), .A1 (n_85), .A2 (a[19]));
NAND2_X1 i_66 (.ZN (n_47), .A1 (n_48), .A2 (n_88));
INV_X1 i_65 (.ZN (p_0[19]), .A (n_47));
NAND3_X1 i_64 (.ZN (n_46), .A1 (n_86), .A2 (n_122), .A3 (n_108));
AOI21_X1 i_63 (.ZN (p_0[18]), .A (n_84), .B1 (n_46), .B2 (a[18]));
OAI21_X1 i_62 (.ZN (n_45), .A (a[17]), .B1 (n_87), .B2 (a[16]));
NAND2_X1 i_61 (.ZN (n_44), .A1 (n_45), .A2 (n_46));
INV_X1 i_60 (.ZN (p_0[17]), .A (n_44));
XNOR2_X1 i_59 (.ZN (n_43), .A (n_87), .B (a[16]));
INV_X1 i_58 (.ZN (p_0[16]), .A (n_43));
NAND2_X1 i_57 (.ZN (n_42), .A1 (n_135), .A2 (n_134));
INV_X1 i_56 (.ZN (n_41), .A (n_42));
NAND2_X1 i_55 (.ZN (n_40), .A1 (n_140), .A2 (n_120));
INV_X1 i_54 (.ZN (n_39), .A (n_40));
NAND2_X1 i_53 (.ZN (n_38), .A1 (n_39), .A2 (n_126));
INV_X1 i_52 (.ZN (n_37), .A (n_38));
NAND4_X1 i_51 (.ZN (n_36), .A1 (n_37), .A2 (n_138), .A3 (n_133), .A4 (n_41));
INV_X1 i_50 (.ZN (n_35), .A (n_36));
INV_X1 i_49 (.ZN (n_34), .A (n_137));
NAND4_X1 i_48 (.ZN (n_33), .A1 (n_37), .A2 (n_133), .A3 (n_34), .A4 (n_41));
OAI21_X1 i_47 (.ZN (n_32), .A (n_33), .B1 (n_35), .B2 (n_139));
INV_X1 i_46 (.ZN (p_0[15]), .A (n_32));
NAND2_X1 i_45 (.ZN (n_31), .A1 (n_37), .A2 (n_133));
INV_X1 i_44 (.ZN (n_30), .A (n_31));
AOI21_X1 i_43 (.ZN (n_29), .A (n_138), .B1 (n_30), .B2 (n_41));
NOR2_X1 i_42 (.ZN (p_0[14]), .A1 (n_29), .A2 (n_35));
NAND3_X1 i_41 (.ZN (n_28), .A1 (n_37), .A2 (n_134), .A3 (n_133));
INV_X1 i_40 (.ZN (n_27), .A (n_28));
OAI22_X1 i_39 (.ZN (n_26), .A1 (n_135), .A2 (n_27), .B1 (n_31), .B2 (n_42));
INV_X1 i_38 (.ZN (p_0[13]), .A (n_26));
NAND2_X1 i_37 (.ZN (n_25), .A1 (n_31), .A2 (a[12]));
NAND2_X1 i_36 (.ZN (n_24), .A1 (n_25), .A2 (n_28));
INV_X1 i_35 (.ZN (p_0[12]), .A (n_24));
NAND2_X1 i_34 (.ZN (n_23), .A1 (n_38), .A2 (a[11]));
NAND2_X1 i_33 (.ZN (n_22), .A1 (n_31), .A2 (n_23));
INV_X1 i_32 (.ZN (p_0[11]), .A (n_22));
NAND3_X1 i_31 (.ZN (n_21), .A1 (n_39), .A2 (n_129), .A3 (n_128));
AOI21_X1 i_30 (.ZN (p_0[10]), .A (n_37), .B1 (n_21), .B2 (a[10]));
NAND2_X1 i_29 (.ZN (n_20), .A1 (n_39), .A2 (n_128));
NAND2_X1 i_28 (.ZN (n_19), .A1 (n_20), .A2 (a[9]));
NAND2_X1 i_27 (.ZN (n_18), .A1 (n_19), .A2 (n_21));
INV_X1 i_26 (.ZN (p_0[9]), .A (n_18));
NAND2_X1 i_25 (.ZN (n_17), .A1 (n_40), .A2 (a[8]));
NAND2_X1 i_24 (.ZN (n_16), .A1 (n_20), .A2 (n_17));
INV_X1 i_23 (.ZN (p_0[8]), .A (n_16));
NOR2_X1 i_22 (.ZN (n_15), .A1 (n_141), .A2 (a[4]));
NAND3_X1 i_21 (.ZN (n_14), .A1 (n_15), .A2 (n_124), .A3 (n_104));
XNOR2_X1 i_20 (.ZN (p_0[7]), .A (n_14), .B (n_125));
INV_X1 i_19 (.ZN (n_13), .A (n_15));
OAI21_X1 i_18 (.ZN (n_12), .A (a[6]), .B1 (n_13), .B2 (a[5]));
NAND2_X1 i_17 (.ZN (n_11), .A1 (n_12), .A2 (n_14));
INV_X1 i_16 (.ZN (p_0[6]), .A (n_11));
XNOR2_X1 i_15 (.ZN (n_10), .A (n_15), .B (n_104));
INV_X1 i_14 (.ZN (p_0[5]), .A (n_10));
NAND2_X1 i_13 (.ZN (n_9), .A1 (n_141), .A2 (a[4]));
NAND2_X1 i_12 (.ZN (n_8), .A1 (n_13), .A2 (n_9));
INV_X1 i_11 (.ZN (p_0[4]), .A (n_8));
NAND3_X1 i_10 (.ZN (n_7), .A1 (n_142), .A2 (n_144), .A3 (n_143));
NAND2_X1 i_9 (.ZN (n_6), .A1 (n_7), .A2 (a[3]));
NAND2_X1 i_8 (.ZN (n_5), .A1 (n_6), .A2 (n_141));
INV_X1 i_7 (.ZN (p_0[3]), .A (n_5));
NAND2_X1 i_6 (.ZN (n_4), .A1 (n_142), .A2 (n_143));
NAND2_X1 i_5 (.ZN (n_3), .A1 (n_4), .A2 (a[2]));
NAND2_X1 i_4 (.ZN (n_2), .A1 (n_3), .A2 (n_7));
INV_X1 i_3 (.ZN (p_0[2]), .A (n_2));
NAND2_X1 i_2 (.ZN (n_1), .A1 (a[0]), .A2 (a[1]));
NAND2_X1 i_1 (.ZN (n_0), .A1 (n_4), .A2 (n_1));
INV_X1 i_0 (.ZN (p_0[1]), .A (n_0));

endmodule //datapath__0_3

module datapath__0_4 (p_0, b);

output [31:0] p_0;
input [31:0] b;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (b[25]));
INV_X1 i_63 (.ZN (n_32), .A (b[21]));
INV_X1 i_62 (.ZN (n_31), .A (b[14]));
INV_X1 i_61 (.ZN (n_30), .A (b[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (b[2]), .A2 (b[1]), .A3 (b[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (b[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (b[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (b[5]), .A3 (b[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (b[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (b[8]), .A3 (b[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (b[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (b[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (b[12]), .A3 (b[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (b[15]), .A3 (b[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (b[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (b[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (b[18]), .A3 (b[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (b[18]), .A3 (b[19]), .A4 (b[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (b[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (b[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (b[23]), .A3 (b[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (b[26]), .A3 (b[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (b[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (b[28]), .A3 (b[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (b[28]), .A3 (b[29]), .A4 (b[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (b[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (b[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (b[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (b[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (b[27]), .B1 (n_9), .B2 (b[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (b[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (b[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (b[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (b[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (b[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (b[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (b[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (b[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (b[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (b[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (b[16]), .B1 (n_19), .B2 (b[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (b[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (b[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (b[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (b[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (b[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (b[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (b[9]), .B1 (n_25), .B2 (b[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (b[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (b[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (b[6]), .B1 (n_27), .B2 (b[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (b[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (b[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (b[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (b[2]), .B1 (b[1]), .B2 (b[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (b[1]), .B (b[0]));

endmodule //datapath__0_4

module halfAdder (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder

module fullAdder (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder

module fullAdder__3_89 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_89

module fullAdder__3_86 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_86

module fullAdder__3_83 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_83

module fullAdder__3_80 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_80

module fullAdder__3_77 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_77

module fullAdder__3_74 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_74

module fullAdder__3_71 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_71

module fullAdder__3_68 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_68

module fullAdder__3_65 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_65

module fullAdder__3_62 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_62

module fullAdder__3_59 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_59

module fullAdder__3_56 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_56

module fullAdder__3_53 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_53

module fullAdder__3_50 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_50

module fullAdder__3_47 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_47

module fullAdder__3_44 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_44

module fullAdder__3_41 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_41

module fullAdder__3_38 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_38

module fullAdder__3_35 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_35

module fullAdder__3_32 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;


XOR2_X1 i_0_3 (.Z (n_0_1), .A (cin), .B (x));
XOR2_X1 i_0_2 (.Z (sum), .A (y), .B (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_32

module fullAdder__3_29 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_29

module fullAdder__3_26 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_26

module fullAdder__3_23 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_23

module fullAdder__3_20 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_20

module fullAdder__3_17 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_17

module fullAdder__3_14 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_14

module fullAdder__3_11 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_11

module fullAdder__3_8 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__3_8

module fullAdder__3_5 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;


OR2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_3), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));

endmodule //fullAdder__3_5

module fullAdder__3_2 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


XOR2_X1 i_0_0 (.Z (sum), .A (cin), .B (y));
AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (cin));

endmodule //fullAdder__3_2

module PartialAdder (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__3_89 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__3_86 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__3_83 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__3_80 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__3_77 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__3_74 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__3_71 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__3_68 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__3_65 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__3_62 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__3_59 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__3_56 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__3_53 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__3_50 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__3_47 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__3_44 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__3_41 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__3_38 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__3_35 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__3_32 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__3_29 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__3_26 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__3_23 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__3_20 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__3_17 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__3_14 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__3_11 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__3_8 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__3_5 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__3_2 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .y (b[31]));

endmodule //PartialAdder

module datapath (b, a, p_0);

output [32:0] p_0;
input [31:0] a;
input [31:0] b;
wire n_0;
wire n_193;
wire n_88;
wire n_124;
wire n_4;
wire n_5;
wire n_9;
wire n_111;
wire n_117;
wire n_6;
wire n_8;
wire n_113;
wire n_110;
wire n_7;
wire n_11;
wire n_112;
wire n_10;
wire n_89;
wire n_90;
wire n_116;
wire n_109;
wire n_12;
wire n_13;
wire n_130;
wire n_20;
wire n_107;
wire n_14;
wire n_18;
wire n_106;
wire n_108;
wire n_17;
wire n_91;
wire n_16;
wire n_94;
wire n_93;
wire n_21;
wire n_105;
wire n_19;
wire n_132;
wire n_131;
wire n_92;
wire n_101;
wire n_137;
wire n_26;
wire n_27;
wire n_28;
wire n_139;
wire n_104;
wire n_102;
wire n_103;
wire n_42;
wire n_41;
wire n_164;
wire n_166;
wire n_165;
wire n_160;
wire n_64;
wire n_65;
wire n_100;
wire n_99;
wire n_192;
wire n_67;
wire n_66;
wire n_182;
wire n_181;
wire n_98;
wire n_69;
wire n_68;
wire n_71;
wire n_73;
wire n_70;
wire n_72;
wire n_204;
wire n_180;
wire n_74;
wire n_77;
wire n_75;
wire n_76;
wire n_79;
wire n_78;
wire n_82;
wire n_207;
wire n_183;
wire n_179;
wire n_208;
wire n_211;
wire n_189;
wire n_203;
wire n_184;
wire n_114;
wire n_154;
wire n_187;
wire n_15;
wire n_22;
wire n_39;
wire n_38;
wire n_51;
wire n_194;
wire n_53;
wire n_195;
wire n_52;
wire n_48;
wire n_196;
wire n_50;
wire n_197;
wire n_45;
wire n_49;
wire n_198;
wire n_47;
wire n_199;
wire n_46;
wire n_40;
wire n_200;
wire n_44;
wire n_201;
wire n_43;
wire n_202;
wire n_37;
wire n_205;
wire n_33;
wire n_206;
wire n_35;
wire n_34;
wire n_210;
wire n_25;
wire n_30;
wire n_1;
wire n_31;
wire n_24;
wire n_23;
wire n_55;
wire n_54;
wire n_29;
wire n_58;
wire n_57;
wire n_36;
wire n_32;
wire n_56;
wire n_60;
wire n_63;
wire n_59;
wire n_62;
wire n_61;
wire n_81;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_97;
wire n_95;
wire n_96;
wire n_115;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_138;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_146;
wire n_145;
wire n_149;
wire n_148;
wire n_147;
wire n_150;
wire n_152;
wire n_151;
wire n_161;
wire n_156;
wire n_153;
wire n_159;
wire n_155;
wire n_158;
wire n_157;
wire n_163;
wire n_162;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_175;
wire n_172;
wire n_174;
wire n_173;
wire n_177;
wire n_176;
wire n_178;
wire n_186;
wire n_185;
wire n_188;
wire n_191;
wire n_190;
wire n_209;


NAND2_X1 i_244 (.ZN (n_211), .A1 (b[31]), .A2 (a[31]));
NOR2_X1 i_243 (.ZN (n_209), .A1 (b[31]), .A2 (a[31]));
INV_X1 i_242 (.ZN (n_208), .A (n_209));
NOR2_X1 i_241 (.ZN (n_207), .A1 (b[30]), .A2 (a[30]));
INV_X1 i_240 (.ZN (n_204), .A (n_207));
NAND3_X1 i_239 (.ZN (n_203), .A1 (n_182), .A2 (n_204), .A3 (n_208));
NAND2_X1 i_238 (.ZN (n_192), .A1 (b[28]), .A2 (a[28]));
AOI21_X1 i_237 (.ZN (n_191), .A (n_203), .B1 (n_181), .B2 (n_192));
OAI21_X1 i_236 (.ZN (n_190), .A (n_211), .B1 (n_180), .B2 (n_209));
NOR2_X1 i_235 (.ZN (n_189), .A1 (n_191), .A2 (n_190));
NAND3_X1 i_234 (.ZN (n_188), .A1 (n_164), .A2 (n_167), .A3 (n_177));
AOI21_X1 i_233 (.ZN (n_187), .A (n_188), .B1 (n_163), .B2 (n_162));
AOI21_X1 i_232 (.ZN (n_186), .A (n_188), .B1 (n_160), .B2 (n_166));
OAI21_X1 i_231 (.ZN (n_185), .A (n_176), .B1 (n_178), .B2 (n_168));
AOI211_X1 i_230 (.ZN (n_184), .A (n_186), .B (n_185), .C1 (n_155), .C2 (n_187));
NOR2_X1 i_229 (.ZN (n_183), .A1 (b[29]), .A2 (a[29]));
INV_X1 i_228 (.ZN (n_182), .A (n_183));
NAND2_X1 i_227 (.ZN (n_181), .A1 (b[29]), .A2 (a[29]));
NAND2_X1 i_226 (.ZN (n_180), .A1 (b[30]), .A2 (a[30]));
AND3_X1 i_225 (.ZN (n_179), .A1 (n_182), .A2 (n_180), .A3 (n_181));
NOR2_X1 i_224 (.ZN (n_178), .A1 (b[27]), .A2 (a[27]));
INV_X1 i_223 (.ZN (n_177), .A (n_178));
NAND2_X1 i_222 (.ZN (n_176), .A1 (b[27]), .A2 (a[27]));
NAND2_X1 i_221 (.ZN (n_175), .A1 (n_177), .A2 (n_176));
NAND2_X1 i_220 (.ZN (n_174), .A1 (n_164), .A2 (n_167));
AND3_X1 i_219 (.ZN (n_173), .A1 (n_165), .A2 (n_160), .A3 (n_166));
OAI21_X1 i_218 (.ZN (n_172), .A (n_168), .B1 (n_174), .B2 (n_173));
XNOR2_X1 i_216 (.ZN (p_0[27]), .A (n_175), .B (n_172));
XOR2_X1 i_215 (.Z (p_0[26]), .A (n_170), .B (n_171));
NAND2_X1 i_214 (.ZN (n_171), .A1 (n_167), .A2 (n_168));
NAND2_X1 i_213 (.ZN (n_170), .A1 (n_169), .A2 (n_164));
NAND3_X1 i_212 (.ZN (n_169), .A1 (n_166), .A2 (n_165), .A3 (n_160));
NAND2_X1 i_211 (.ZN (n_168), .A1 (a[26]), .A2 (b[26]));
OR2_X1 i_210 (.ZN (n_167), .A1 (a[26]), .A2 (b[26]));
NAND2_X1 i_209 (.ZN (n_166), .A1 (a[25]), .A2 (b[25]));
NAND2_X1 i_208 (.ZN (n_165), .A1 (n_152), .A2 (n_161));
OR2_X1 i_207 (.ZN (n_164), .A1 (a[25]), .A2 (b[25]));
INV_X1 i_206 (.ZN (n_163), .A (b[24]));
INV_X1 i_205 (.ZN (n_162), .A (a[24]));
NAND2_X1 i_204 (.ZN (n_161), .A1 (n_163), .A2 (n_162));
NAND2_X1 i_203 (.ZN (n_160), .A1 (b[24]), .A2 (a[24]));
NAND3_X1 i_202 (.ZN (n_159), .A1 (n_139), .A2 (n_142), .A3 (n_149));
AOI21_X1 i_201 (.ZN (n_158), .A (n_159), .B1 (n_102), .B2 (n_104));
OAI21_X1 i_200 (.ZN (n_157), .A (n_148), .B1 (n_150), .B2 (n_143));
NOR2_X1 i_199 (.ZN (n_156), .A1 (n_158), .A2 (n_157));
INV_X1 i_198 (.ZN (n_155), .A (n_156));
NOR2_X1 i_197 (.ZN (n_154), .A1 (n_103), .A2 (n_159));
INV_X1 i_196 (.ZN (n_153), .A (n_154));
OAI21_X1 i_195 (.ZN (n_152), .A (n_156), .B1 (n_137), .B2 (n_153));
NAND2_X1 i_194 (.ZN (n_151), .A1 (n_161), .A2 (n_160));
XNOR2_X1 i_193 (.ZN (p_0[24]), .A (n_152), .B (n_151));
NOR2_X1 i_192 (.ZN (n_150), .A1 (a[23]), .A2 (b[23]));
INV_X1 i_191 (.ZN (n_149), .A (n_150));
NAND2_X1 i_190 (.ZN (n_148), .A1 (a[23]), .A2 (b[23]));
NAND2_X1 i_189 (.ZN (n_147), .A1 (n_138), .A2 (n_139));
AOI21_X1 i_188 (.ZN (n_146), .A (n_140), .B1 (n_143), .B2 (n_147));
NAND2_X1 i_187 (.ZN (n_145), .A1 (n_149), .A2 (n_148));
XNOR2_X2 i_186 (.ZN (p_0[23]), .A (n_146), .B (n_145));
XOR2_X1 i_185 (.Z (p_0[22]), .A (n_141), .B (n_144));
NAND2_X1 i_184 (.ZN (n_144), .A1 (n_142), .A2 (n_143));
NAND2_X1 i_183 (.ZN (n_143), .A1 (a[22]), .A2 (b[22]));
INV_X1 i_182 (.ZN (n_142), .A (n_140));
NAND2_X1 i_181 (.ZN (n_141), .A1 (n_138), .A2 (n_139));
NOR2_X1 i_180 (.ZN (n_140), .A1 (a[22]), .A2 (b[22]));
OR2_X1 i_179 (.ZN (n_139), .A1 (a[21]), .A2 (b[21]));
OAI211_X2 i_178 (.ZN (n_138), .A (n_102), .B (n_104), .C1 (n_137), .C2 (n_103));
AOI211_X2 i_177 (.ZN (n_137), .A (n_134), .B (n_135), .C1 (n_130), .C2 (n_136));
AOI21_X1 i_176 (.ZN (n_136), .A (n_133), .B1 (n_131), .B2 (n_132));
OAI21_X1 i_175 (.ZN (n_135), .A (n_95), .B1 (n_97), .B2 (n_92));
AOI21_X1 i_174 (.ZN (n_134), .A (n_133), .B1 (n_107), .B2 (n_108));
NAND3_X1 i_173 (.ZN (n_133), .A1 (n_106), .A2 (n_96), .A3 (n_93));
INV_X1 i_172 (.ZN (n_132), .A (b[16]));
INV_X1 i_171 (.ZN (n_131), .A (a[16]));
OR4_X2 i_170 (.ZN (n_130), .A1 (n_126), .A2 (n_127), .A3 (n_128), .A4 (n_129));
AOI21_X1 i_169 (.ZN (n_129), .A (n_125), .B1 (n_89), .B2 (n_117));
NOR2_X1 i_168 (.ZN (n_128), .A1 (n_110), .A2 (n_115));
INV_X1 i_167 (.ZN (n_127), .A (n_109));
NOR3_X1 i_166 (.ZN (n_126), .A1 (n_124), .A2 (n_90), .A3 (n_125));
NAND3_X1 i_165 (.ZN (n_125), .A1 (n_116), .A2 (n_111), .A3 (n_113));
NOR4_X2 i_164 (.ZN (n_124), .A1 (n_120), .A2 (n_121), .A3 (n_122), .A4 (n_123));
NOR2_X1 i_163 (.ZN (n_123), .A1 (n_81), .A2 (n_62));
INV_X1 i_162 (.ZN (n_122), .A (n_84));
AOI21_X1 i_161 (.ZN (n_121), .A (n_119), .B1 (n_25), .B2 (n_54));
AOI211_X1 i_160 (.ZN (n_120), .A (n_118), .B (n_119), .C1 (n_57), .C2 (n_58));
NAND3_X1 i_159 (.ZN (n_119), .A1 (n_55), .A2 (n_83), .A3 (n_61));
INV_X2 i_158 (.ZN (n_118), .A (n_31));
NAND2_X1 i_157 (.ZN (n_117), .A1 (a[13]), .A2 (b[13]));
INV_X1 i_156 (.ZN (n_116), .A (n_115));
NOR2_X1 i_155 (.ZN (n_115), .A1 (a[15]), .A2 (b[15]));
INV_X1 i_154 (.ZN (n_113), .A (n_112));
NOR2_X1 i_153 (.ZN (n_112), .A1 (a[14]), .A2 (b[14]));
OR2_X1 i_152 (.ZN (n_111), .A1 (a[13]), .A2 (b[13]));
NAND2_X1 i_151 (.ZN (n_110), .A1 (a[14]), .A2 (b[14]));
NAND2_X1 i_150 (.ZN (n_109), .A1 (a[15]), .A2 (b[15]));
NAND2_X1 i_149 (.ZN (n_108), .A1 (a[17]), .A2 (b[17]));
NAND2_X1 i_148 (.ZN (n_107), .A1 (a[16]), .A2 (b[16]));
INV_X1 i_147 (.ZN (n_106), .A (n_105));
NOR2_X1 i_146 (.ZN (n_105), .A1 (a[17]), .A2 (b[17]));
NAND2_X1 i_145 (.ZN (n_104), .A1 (a[21]), .A2 (b[21]));
NOR2_X1 i_144 (.ZN (n_103), .A1 (a[20]), .A2 (b[20]));
NAND2_X1 i_143 (.ZN (n_102), .A1 (a[20]), .A2 (b[20]));
OAI21_X1 i_142 (.ZN (n_101), .A (n_102), .B1 (a[20]), .B2 (b[20]));
NOR2_X1 i_141 (.ZN (n_97), .A1 (a[19]), .A2 (b[19]));
INV_X1 i_140 (.ZN (n_96), .A (n_97));
NAND2_X1 i_139 (.ZN (n_95), .A1 (a[19]), .A2 (b[19]));
AOI21_X1 i_138 (.ZN (n_94), .A (n_97), .B1 (a[19]), .B2 (b[19]));
OR2_X1 i_137 (.ZN (n_93), .A1 (a[18]), .A2 (b[18]));
NAND2_X1 i_136 (.ZN (n_92), .A1 (a[18]), .A2 (b[18]));
NAND2_X1 i_135 (.ZN (n_91), .A1 (n_93), .A2 (n_92));
NOR2_X1 i_134 (.ZN (n_90), .A1 (b[12]), .A2 (a[12]));
NAND2_X1 i_133 (.ZN (n_89), .A1 (b[12]), .A2 (a[12]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_89), .B1 (b[12]), .B2 (a[12]));
XNOR2_X1 i_131 (.ZN (p_0[11]), .A (n_86), .B (n_87));
NAND2_X1 i_130 (.ZN (n_87), .A1 (n_83), .A2 (n_84));
NAND2_X1 i_129 (.ZN (n_86), .A1 (n_85), .A2 (n_62));
NAND3_X1 i_128 (.ZN (n_85), .A1 (n_61), .A2 (n_55), .A3 (n_63));
NAND2_X1 i_127 (.ZN (n_84), .A1 (a[11]), .A2 (b[11]));
INV_X1 i_126 (.ZN (n_83), .A (n_81));
NOR2_X1 i_125 (.ZN (n_81), .A1 (a[11]), .A2 (b[11]));
NAND3_X1 i_123 (.ZN (n_63), .A1 (n_29), .A2 (n_54), .A3 (n_25));
NAND2_X1 i_122 (.ZN (n_62), .A1 (a[10]), .A2 (b[10]));
OR2_X1 i_121 (.ZN (n_61), .A1 (a[10]), .A2 (b[10]));
AOI22_X1 i_120 (.ZN (n_60), .A1 (n_62), .A2 (n_61), .B1 (n_55), .B2 (n_24));
AND3_X1 i_119 (.ZN (n_59), .A1 (n_62), .A2 (n_61), .A3 (n_55));
AOI22_X1 i_118 (.ZN (p_0[10]), .A1 (n_54), .A2 (n_60), .B1 (n_63), .B2 (n_59));
INV_X1 i_117 (.ZN (n_58), .A (b[8]));
INV_X1 i_116 (.ZN (n_57), .A (a[8]));
NOR2_X1 i_115 (.ZN (n_56), .A1 (b[9]), .A2 (a[9]));
INV_X1 i_114 (.ZN (n_55), .A (n_56));
NAND2_X1 i_113 (.ZN (n_54), .A1 (b[9]), .A2 (a[9]));
NAND2_X2 i_112 (.ZN (n_53), .A1 (n_15), .A2 (n_22));
OR2_X1 i_111 (.ZN (n_52), .A1 (b[2]), .A2 (a[2]));
OR2_X2 i_110 (.ZN (n_51), .A1 (b[1]), .A2 (a[1]));
NAND3_X2 i_109 (.ZN (n_50), .A1 (n_53), .A2 (n_51), .A3 (n_52));
NAND2_X1 i_108 (.ZN (n_49), .A1 (b[3]), .A2 (a[3]));
NAND2_X1 i_107 (.ZN (n_48), .A1 (b[2]), .A2 (a[2]));
NAND3_X2 i_106 (.ZN (n_47), .A1 (n_50), .A2 (n_49), .A3 (n_48));
OR2_X1 i_105 (.ZN (n_46), .A1 (b[4]), .A2 (a[4]));
OR2_X1 i_104 (.ZN (n_45), .A1 (b[3]), .A2 (a[3]));
NAND3_X2 i_103 (.ZN (n_44), .A1 (n_47), .A2 (n_46), .A3 (n_45));
NAND2_X1 i_102 (.ZN (n_43), .A1 (b[5]), .A2 (a[5]));
NAND2_X1 i_101 (.ZN (n_40), .A1 (b[4]), .A2 (a[4]));
NAND3_X2 i_100 (.ZN (n_39), .A1 (n_44), .A2 (n_43), .A3 (n_40));
OR2_X1 i_99 (.ZN (n_38), .A1 (b[5]), .A2 (a[5]));
OR2_X1 i_98 (.ZN (n_37), .A1 (b[6]), .A2 (a[6]));
NOR2_X1 i_97 (.ZN (n_36), .A1 (b[7]), .A2 (a[7]));
INV_X1 i_96 (.ZN (n_35), .A (n_36));
NAND2_X1 i_95 (.ZN (n_34), .A1 (b[7]), .A2 (a[7]));
NAND2_X1 i_94 (.ZN (n_33), .A1 (b[6]), .A2 (a[6]));
NAND3_X1 i_93 (.ZN (n_32), .A1 (n_39), .A2 (n_38), .A3 (n_37));
OAI221_X2 i_92 (.ZN (n_31), .A (n_34), .B1 (n_36), .B2 (n_33), .C1 (n_36), .C2 (n_32));
NAND2_X1 i_91 (.ZN (n_30), .A1 (n_58), .A2 (n_57));
NAND2_X1 i_90 (.ZN (n_29), .A1 (n_31), .A2 (n_30));
NAND2_X1 i_89 (.ZN (n_25), .A1 (b[8]), .A2 (a[8]));
NAND2_X1 i_88 (.ZN (n_24), .A1 (n_29), .A2 (n_25));
NAND2_X1 i_87 (.ZN (n_23), .A1 (n_55), .A2 (n_54));
XNOR2_X1 i_86 (.ZN (p_0[9]), .A (n_24), .B (n_23));
XNOR2_X1 i_83 (.ZN (p_0[8]), .A (n_31), .B (n_1));
NAND2_X1 i_82 (.ZN (n_1), .A1 (n_25), .A2 (n_30));
XNOR2_X1 i_81 (.ZN (p_0[7]), .A (n_206), .B (n_210));
NAND2_X1 i_80 (.ZN (n_210), .A1 (n_35), .A2 (n_34));
NAND2_X1 i_79 (.ZN (n_206), .A1 (n_205), .A2 (n_33));
NAND3_X1 i_78 (.ZN (n_205), .A1 (n_39), .A2 (n_38), .A3 (n_37));
XNOR2_X1 i_77 (.ZN (p_0[5]), .A (n_201), .B (n_202));
NAND2_X1 i_76 (.ZN (n_202), .A1 (n_38), .A2 (n_43));
NAND2_X1 i_75 (.ZN (n_201), .A1 (n_44), .A2 (n_40));
XOR2_X1 i_74 (.Z (p_0[4]), .A (n_199), .B (n_200));
NAND2_X1 i_73 (.ZN (n_200), .A1 (n_46), .A2 (n_40));
NAND2_X1 i_72 (.ZN (n_199), .A1 (n_47), .A2 (n_45));
XNOR2_X1 i_71 (.ZN (p_0[3]), .A (n_197), .B (n_198));
NAND2_X1 i_70 (.ZN (n_198), .A1 (n_45), .A2 (n_49));
NAND2_X1 i_69 (.ZN (n_197), .A1 (n_50), .A2 (n_48));
XOR2_X1 i_68 (.Z (p_0[2]), .A (n_195), .B (n_196));
NAND2_X1 i_67 (.ZN (n_196), .A1 (n_52), .A2 (n_48));
NAND2_X1 i_66 (.ZN (n_195), .A1 (n_53), .A2 (n_51));
XOR2_X1 i_65 (.Z (p_0[1]), .A (n_194), .B (n_15));
NAND2_X1 i_64 (.ZN (n_194), .A1 (n_51), .A2 (n_22));
XOR2_X1 i_217 (.Z (p_0[0]), .A (b[0]), .B (a[0]));
NAND2_X1 i_63 (.ZN (n_193), .A1 (n_39), .A2 (n_38));
NAND2_X1 i_62 (.ZN (n_22), .A1 (b[1]), .A2 (a[1]));
NAND2_X2 i_61 (.ZN (n_15), .A1 (b[0]), .A2 (a[0]));
NAND2_X1 i_60 (.ZN (n_114), .A1 (n_154), .A2 (n_187));
OAI21_X1 i_59 (.ZN (n_100), .A (n_184), .B1 (n_137), .B2 (n_114));
OR2_X1 i_58 (.ZN (n_99), .A1 (a[28]), .A2 (b[28]));
NAND2_X1 i_57 (.ZN (n_98), .A1 (n_100), .A2 (n_99));
OAI21_X1 i_56 (.ZN (p_0[32]), .A (n_189), .B1 (n_98), .B2 (n_203));
NAND2_X1 i_55 (.ZN (n_82), .A1 (n_208), .A2 (n_211));
NAND3_X1 i_54 (.ZN (n_79), .A1 (n_98), .A2 (n_192), .A3 (n_179));
AOI21_X1 i_53 (.ZN (n_78), .A (n_207), .B1 (n_183), .B2 (n_180));
NAND3_X1 i_52 (.ZN (n_77), .A1 (n_79), .A2 (n_82), .A3 (n_78));
INV_X1 i_51 (.ZN (n_76), .A (n_82));
NAND2_X1 i_50 (.ZN (n_75), .A1 (n_79), .A2 (n_78));
NAND2_X1 i_49 (.ZN (n_74), .A1 (n_75), .A2 (n_76));
NAND2_X1 i_48 (.ZN (p_0[31]), .A1 (n_74), .A2 (n_77));
NAND2_X1 i_47 (.ZN (n_73), .A1 (n_204), .A2 (n_180));
INV_X1 i_46 (.ZN (n_72), .A (n_73));
NAND3_X1 i_45 (.ZN (n_71), .A1 (n_98), .A2 (n_192), .A3 (n_181));
NAND2_X1 i_44 (.ZN (n_70), .A1 (n_71), .A2 (n_182));
NAND2_X1 i_43 (.ZN (n_69), .A1 (n_70), .A2 (n_72));
NAND3_X1 i_42 (.ZN (n_68), .A1 (n_71), .A2 (n_182), .A3 (n_73));
NAND2_X1 i_41 (.ZN (p_0[30]), .A1 (n_69), .A2 (n_68));
NAND2_X1 i_40 (.ZN (n_67), .A1 (n_98), .A2 (n_192));
NAND2_X1 i_39 (.ZN (n_66), .A1 (n_182), .A2 (n_181));
XNOR2_X1 i_38 (.ZN (p_0[29]), .A (n_67), .B (n_66));
NAND2_X1 i_37 (.ZN (n_65), .A1 (n_99), .A2 (n_192));
XOR2_X1 i_36 (.Z (n_64), .A (n_65), .B (n_100));
INV_X1 i_35 (.ZN (p_0[28]), .A (n_64));
NAND2_X1 i_34 (.ZN (n_42), .A1 (n_165), .A2 (n_160));
NAND2_X1 i_33 (.ZN (n_41), .A1 (n_164), .A2 (n_166));
XNOR2_X1 i_32 (.ZN (p_0[25]), .A (n_42), .B (n_41));
OAI21_X1 i_31 (.ZN (n_28), .A (n_102), .B1 (n_137), .B2 (n_103));
NAND2_X1 i_30 (.ZN (n_27), .A1 (n_139), .A2 (n_104));
XOR2_X1 i_29 (.Z (n_26), .A (n_27), .B (n_28));
INV_X1 i_28 (.ZN (p_0[21]), .A (n_26));
XOR2_X1 i_27 (.Z (p_0[20]), .A (n_101), .B (n_137));
INV_X1 i_26 (.ZN (n_21), .A (n_92));
NAND2_X1 i_25 (.ZN (n_20), .A1 (n_132), .A2 (n_131));
INV_X1 i_24 (.ZN (n_19), .A (n_107));
AOI21_X1 i_23 (.ZN (n_18), .A (n_19), .B1 (n_130), .B2 (n_20));
AOI21_X1 i_22 (.ZN (n_17), .A (n_105), .B1 (n_18), .B2 (n_108));
OAI21_X1 i_21 (.ZN (n_16), .A (n_93), .B1 (n_17), .B2 (n_21));
XNOR2_X1 i_20 (.ZN (p_0[19]), .A (n_16), .B (n_94));
XNOR2_X1 i_19 (.ZN (p_0[18]), .A (n_17), .B (n_91));
NAND2_X1 i_18 (.ZN (n_14), .A1 (n_106), .A2 (n_108));
XOR2_X1 i_17 (.Z (p_0[17]), .A (n_14), .B (n_18));
NAND2_X1 i_16 (.ZN (n_13), .A1 (n_20), .A2 (n_107));
XOR2_X1 i_15 (.Z (n_12), .A (n_13), .B (n_130));
INV_X1 i_14 (.ZN (p_0[16]), .A (n_12));
NAND2_X1 i_13 (.ZN (n_11), .A1 (n_116), .A2 (n_109));
INV_X1 i_12 (.ZN (n_10), .A (n_117));
OAI21_X1 i_11 (.ZN (n_9), .A (n_89), .B1 (n_124), .B2 (n_90));
OAI21_X1 i_10 (.ZN (n_8), .A (n_111), .B1 (n_9), .B2 (n_10));
AOI21_X1 i_9 (.ZN (n_7), .A (n_112), .B1 (n_8), .B2 (n_110));
XNOR2_X1 i_8 (.ZN (p_0[15]), .A (n_7), .B (n_11));
NAND2_X1 i_7 (.ZN (n_6), .A1 (n_113), .A2 (n_110));
XOR2_X1 i_6 (.Z (p_0[14]), .A (n_6), .B (n_8));
NAND2_X1 i_5 (.ZN (n_5), .A1 (n_111), .A2 (n_117));
XOR2_X1 i_4 (.Z (n_4), .A (n_5), .B (n_9));
INV_X1 i_3 (.ZN (p_0[13]), .A (n_4));
XOR2_X1 i_2 (.Z (p_0[12]), .A (n_88), .B (n_124));
NAND2_X1 i_1 (.ZN (n_0), .A1 (n_37), .A2 (n_33));
XOR2_X1 i_0 (.Z (p_0[6]), .A (n_0), .B (n_193));

endmodule //datapath

module adderPlus (a, b, sum, cout);

output cout;
output [31:0] sum;
input [31:0] a;
input [31:0] b;


datapath i_0 (.p_0 ({cout, sum[31], sum[30], sum[29], sum[28], sum[27], sum[26], 
    sum[25], sum[24], sum[23], sum[22], sum[21], sum[20], sum[19], sum[18], sum[17], 
    sum[16], sum[15], sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
    sum[7], sum[6], sum[5], sum[4], sum[3], sum[2], sum[1], sum[0]}), .a ({a[31], 
    a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], a[21], a[20], 
    a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8], 
    a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), .b ({b[31], b[30], b[29], b[28], 
    b[27], b[26], b[25], b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], 
    b[16], b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], 
    b[4], b[3], b[2], b[1], b[0]}));

endmodule //adderPlus

module halfAdder__0_43 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X2 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__0_43

module fullAdder__0_46 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__0_46

module fullAdder__1_89 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (y), .A2 (cin));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (x), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (x), .A3 (n_0_5));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_3 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_4));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_7), .B2 (n_0_1));

endmodule //fullAdder__1_89

module fullAdder__1_86 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


OAI21_X1 i_0_8 (.ZN (sum), .A (n_0_5), .B1 (n_0_6), .B2 (y));
AND2_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_3), .A2 (n_0_4));
NAND3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1));
OR2_X1 i_0_3 (.ZN (n_0_3), .A1 (x), .A2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_86

module fullAdder__1_83 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_5), .B2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_4));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_83

module fullAdder__1_80 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
XNOR2_X1 i_0_7 (.ZN (n_0_5), .A (y), .B (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_80

module fullAdder__1_77 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_77

module fullAdder__1_74 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_3), .B1 (x), .B2 (n_0_2));
INV_X1 i_0_5 (.ZN (n_0_4), .A (x));
XNOR2_X1 i_0_4 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_3 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_74

module fullAdder__1_71 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (x));
INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_11), .A2 (n_0_9), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_9));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (n_0_10));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (x), .B1 (n_0_5), .B2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_71

module fullAdder__1_68 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_68

module fullAdder__1_65 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_65

module fullAdder__1_62 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_62

module fullAdder__1_59 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_59

module fullAdder__1_56 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_56

module fullAdder__1_53 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_53

module fullAdder__1_50 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_50

module fullAdder__1_47 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_47

module fullAdder__1_44 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_44

module fullAdder__1_41 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_41

module fullAdder__1_38 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_38

module fullAdder__1_35 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_35

module fullAdder__1_32 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_32

module fullAdder__1_29 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_29

module fullAdder__1_26 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_26

module fullAdder__1_23 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_23

module fullAdder__1_20 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_20

module fullAdder__1_17 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_17

module fullAdder__1_14 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_14

module fullAdder__1_11 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_11

module fullAdder__1_8 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_8

module fullAdder__1_5 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_5

module fullAdder__1_2 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2

module PartialAdder__0_47 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__0_43 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__0_46 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_89 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_86 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_83 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_80 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_77 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_74 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_71 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_68 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_65 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_62 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_59 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_56 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_53 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_50 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_47 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_44 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_41 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_38 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_35 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_32 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_29 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_26 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_23 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_20 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_17 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_14 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_11 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_8 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_5 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__0_47

module halfAdder__1_2711 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2711

module fullAdder__1_2714 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2714

module fullAdder__1_2717 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2717

module fullAdder__1_2720 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (x), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (x), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OR2_X1 i_0_4 (.ZN (n_0_3), .A1 (y), .A2 (cin));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));

endmodule //fullAdder__1_2720

module fullAdder__1_2723 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2723

module fullAdder__1_2726 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2726

module fullAdder__1_2729 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2729

module fullAdder__1_2732 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2732

module fullAdder__1_2735 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (x));
INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_11), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2735

module fullAdder__1_2738 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2738

module fullAdder__1_2741 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2741

module fullAdder__1_2744 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2744

module fullAdder__1_2747 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2747

module fullAdder__1_2750 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2750

module fullAdder__1_2753 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2753

module fullAdder__1_2756 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2756

module fullAdder__1_2759 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2759

module fullAdder__1_2762 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2762

module fullAdder__1_2765 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2765

module fullAdder__1_2768 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2768

module fullAdder__1_2771 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2771

module fullAdder__1_2774 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2774

module fullAdder__1_2777 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2777

module fullAdder__1_2780 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2780

module fullAdder__1_2783 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2783

module fullAdder__1_2786 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2786

module fullAdder__1_2789 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2789

module fullAdder__1_2792 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2792

module fullAdder__1_2795 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2795

module fullAdder__1_2798 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2798

module fullAdder__1_2801 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2801

module fullAdder__1_2804 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2804

module PartialAdder__1_2805 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2711 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2714 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2717 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2720 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2723 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2726 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2729 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2732 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2735 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2738 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2741 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2744 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2747 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2750 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2753 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2756 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2759 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2762 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2765 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2768 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2771 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2774 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2777 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2780 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2783 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2786 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2789 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2792 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2795 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2798 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2801 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2804 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2805

module halfAdder__1_2614 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2614

module fullAdder__1_2617 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2617

module fullAdder__1_2620 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_0), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
AOI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (y));
NOR2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_2620

module fullAdder__1_2623 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2623

module fullAdder__1_2626 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2626

module fullAdder__1_2629 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


NAND2_X1 i_0_13 (.ZN (n_0_11), .A1 (y), .A2 (cin));
INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_10), .A2 (n_0_9));
NAND3_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (x), .A3 (n_0_11));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_11));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (n_0_6), .B1 (n_0_5), .B2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_7));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2629

module fullAdder__1_2632 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2632

module fullAdder__1_2635 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2635

module fullAdder__1_2638 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2638

module fullAdder__1_2641 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2641

module fullAdder__1_2644 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2644

module fullAdder__1_2647 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2647

module fullAdder__1_2650 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2650

module fullAdder__1_2653 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2653

module fullAdder__1_2656 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2656

module fullAdder__1_2659 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2659

module fullAdder__1_2662 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2662

module fullAdder__1_2665 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2665

module fullAdder__1_2668 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2668

module fullAdder__1_2671 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2671

module fullAdder__1_2674 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2674

module fullAdder__1_2677 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2677

module fullAdder__1_2680 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2680

module fullAdder__1_2683 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2683

module fullAdder__1_2686 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2686

module fullAdder__1_2689 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2689

module fullAdder__1_2692 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2692

module fullAdder__1_2695 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2695

module fullAdder__1_2698 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2698

module fullAdder__1_2701 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2701

module fullAdder__1_2704 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2704

module fullAdder__1_2707 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2707

module PartialAdder__1_2708 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2614 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2617 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2620 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2623 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2626 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2629 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2632 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2635 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2638 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2641 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2644 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2647 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2650 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2653 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2656 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2659 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2662 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2665 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2668 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2671 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2674 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2677 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2680 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2683 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2686 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2689 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2692 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2695 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2698 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2701 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2704 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2707 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2708

module halfAdder__1_2517 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2517

module fullAdder__1_2520 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X2 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_2520

module fullAdder__1_2523 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2523

module fullAdder__1_2526 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


AOI21_X2 i_0_8 (.ZN (sum), .A (n_0_5), .B1 (n_0_6), .B2 (x));
OR2_X2 i_0_7 (.ZN (n_0_6), .A1 (n_0_3), .A2 (n_0_4));
NOR3_X2 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (x), .A3 (n_0_4));
NOR2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (n_0_2));
AND2_X1 i_0_4 (.ZN (n_0_3), .A1 (y), .A2 (n_0_2));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (x));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_2526

module fullAdder__1_2529 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2529

module fullAdder__1_2532 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_2532

module fullAdder__1_2535 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2535

module fullAdder__1_2538 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2538

module fullAdder__1_2541 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2541

module fullAdder__1_2544 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2544

module fullAdder__1_2547 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2547

module fullAdder__1_2550 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2550

module fullAdder__1_2553 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2553

module fullAdder__1_2556 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2556

module fullAdder__1_2559 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2559

module fullAdder__1_2562 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2562

module fullAdder__1_2565 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2565

module fullAdder__1_2568 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2568

module fullAdder__1_2571 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2571

module fullAdder__1_2574 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2574

module fullAdder__1_2577 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2577

module fullAdder__1_2580 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2580

module fullAdder__1_2583 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2583

module fullAdder__1_2586 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2586

module fullAdder__1_2589 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2589

module fullAdder__1_2592 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2592

module fullAdder__1_2595 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2595

module fullAdder__1_2598 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2598

module fullAdder__1_2601 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2601

module fullAdder__1_2604 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2604

module fullAdder__1_2607 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2607

module fullAdder__1_2610 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2610

module PartialAdder__1_2611 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2517 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2520 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2523 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2526 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2529 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2532 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2535 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2538 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2541 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2544 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2547 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2550 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2553 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2556 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2559 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2562 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2565 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2568 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2571 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2574 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2577 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2580 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2583 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2586 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2589 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2592 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2595 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2598 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2601 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2604 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2607 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2610 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2611

module halfAdder__1_2420 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2420

module fullAdder__1_2423 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2423

module fullAdder__1_2426 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_2426

module fullAdder__1_2429 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;


OAI21_X1 i_0_4 (.ZN (n_0_2), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_2429

module fullAdder__1_2432 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_2432

module fullAdder__1_2435 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2435

module fullAdder__1_2438 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2438

module fullAdder__1_2441 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2441

module fullAdder__1_2444 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2444

module fullAdder__1_2447 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2447

module fullAdder__1_2450 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2450

module fullAdder__1_2453 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2453

module fullAdder__1_2456 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2456

module fullAdder__1_2459 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2459

module fullAdder__1_2462 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2462

module fullAdder__1_2465 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2465

module fullAdder__1_2468 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2468

module fullAdder__1_2471 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2471

module fullAdder__1_2474 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2474

module fullAdder__1_2477 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2477

module fullAdder__1_2480 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2480

module fullAdder__1_2483 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2483

module fullAdder__1_2486 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2486

module fullAdder__1_2489 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2489

module fullAdder__1_2492 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2492

module fullAdder__1_2495 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2495

module fullAdder__1_2498 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2498

module fullAdder__1_2501 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2501

module fullAdder__1_2504 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2504

module fullAdder__1_2507 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2507

module fullAdder__1_2510 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2510

module fullAdder__1_2513 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2513

module PartialAdder__1_2514 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2420 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2423 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2426 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2429 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2432 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2435 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2438 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2441 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2444 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2447 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2450 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2453 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2456 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2459 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2462 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2465 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2468 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2471 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2474 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2477 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2480 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2483 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2486 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2489 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2492 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2495 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2498 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2501 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2504 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2507 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2510 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2513 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2514

module halfAdder__1_2323 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2323

module fullAdder__1_2326 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2326

module fullAdder__1_2329 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2329

module fullAdder__1_2332 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_2332

module fullAdder__1_2335 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2335

module fullAdder__1_2338 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2338

module fullAdder__1_2341 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2341

module fullAdder__1_2344 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2344

module fullAdder__1_2347 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_10), .A2 (n_0_7), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2347

module fullAdder__1_2350 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2350

module fullAdder__1_2353 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2353

module fullAdder__1_2356 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2356

module fullAdder__1_2359 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2359

module fullAdder__1_2362 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2362

module fullAdder__1_2365 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2365

module fullAdder__1_2368 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2368

module fullAdder__1_2371 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2371

module fullAdder__1_2374 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2374

module fullAdder__1_2377 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2377

module fullAdder__1_2380 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2380

module fullAdder__1_2383 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2383

module fullAdder__1_2386 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2386

module fullAdder__1_2389 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2389

module fullAdder__1_2392 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2392

module fullAdder__1_2395 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2395

module fullAdder__1_2398 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2398

module fullAdder__1_2401 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2401

module fullAdder__1_2404 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2404

module fullAdder__1_2407 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2407

module fullAdder__1_2410 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2410

module fullAdder__1_2413 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2413

module fullAdder__1_2416 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2416

module PartialAdder__1_2417 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2323 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2326 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2329 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2332 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2335 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2338 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2341 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2344 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2347 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2350 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2353 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2356 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2359 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2362 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2365 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2368 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2371 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2374 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2377 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2380 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2383 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2386 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2389 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2392 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2395 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2398 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2401 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2404 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2407 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2410 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2413 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2416 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2417

module halfAdder__1_2226 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2226

module fullAdder__1_2229 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2229

module fullAdder__1_2232 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2232

module fullAdder__1_2235 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2235

module fullAdder__1_2238 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2238

module fullAdder__1_2241 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (y), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (y));
INV_X1 i_0_5 (.ZN (n_0_3), .A (cin));
INV_X1 i_0_4 (.ZN (n_0_2), .A (x));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_3));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_4), .A2 (n_0_8), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_5));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_6), .B1 (n_0_4), .B2 (n_0_8));

endmodule //fullAdder__1_2241

module fullAdder__1_2244 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2244

module fullAdder__1_2247 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_6), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_2), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_6));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_2247

module fullAdder__1_2250 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2250

module fullAdder__1_2253 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2253

module fullAdder__1_2256 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2256

module fullAdder__1_2259 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2259

module fullAdder__1_2262 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2262

module fullAdder__1_2265 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2265

module fullAdder__1_2268 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2268

module fullAdder__1_2271 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2271

module fullAdder__1_2274 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2274

module fullAdder__1_2277 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2277

module fullAdder__1_2280 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2280

module fullAdder__1_2283 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2283

module fullAdder__1_2286 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2286

module fullAdder__1_2289 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2289

module fullAdder__1_2292 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2292

module fullAdder__1_2295 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2295

module fullAdder__1_2298 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2298

module fullAdder__1_2301 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2301

module fullAdder__1_2304 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2304

module fullAdder__1_2307 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2307

module fullAdder__1_2310 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2310

module fullAdder__1_2313 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2313

module fullAdder__1_2316 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2316

module fullAdder__1_2319 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2319

module PartialAdder__1_2320 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2226 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2229 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2232 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2235 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2238 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2241 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2244 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2247 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2250 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2253 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2256 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2259 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2262 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2265 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2268 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2271 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2274 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2277 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2280 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2283 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2286 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2289 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2292 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2295 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2298 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2301 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2304 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2307 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2310 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2313 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2316 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2319 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2320

module halfAdder__1_2129 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2129

module fullAdder__1_2132 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


AOI21_X1 i_0_8 (.ZN (sum), .A (n_0_5), .B1 (n_0_6), .B2 (x));
OR2_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_3), .A2 (n_0_4));
NOR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (x), .A3 (n_0_4));
NOR2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (n_0_1));
AND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2132

module fullAdder__1_2135 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2135

module fullAdder__1_2138 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2138

module fullAdder__1_2141 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (x));
INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_11), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_2141

module fullAdder__1_2144 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2144

module fullAdder__1_2147 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2147

module fullAdder__1_2150 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2150

module fullAdder__1_2153 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2153

module fullAdder__1_2156 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (n_0_4), .A3 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_3));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_5), .B1 (n_0_6), .B2 (n_0_3));

endmodule //fullAdder__1_2156

module fullAdder__1_2159 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2159

module fullAdder__1_2162 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2162

module fullAdder__1_2165 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2165

module fullAdder__1_2168 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2168

module fullAdder__1_2171 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2171

module fullAdder__1_2174 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2174

module fullAdder__1_2177 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2177

module fullAdder__1_2180 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2180

module fullAdder__1_2183 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2183

module fullAdder__1_2186 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2186

module fullAdder__1_2189 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2189

module fullAdder__1_2192 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2192

module fullAdder__1_2195 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2195

module fullAdder__1_2198 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2198

module fullAdder__1_2201 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2201

module fullAdder__1_2204 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2204

module fullAdder__1_2207 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2207

module fullAdder__1_2210 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2210

module fullAdder__1_2213 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2213

module fullAdder__1_2216 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2216

module fullAdder__1_2219 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2219

module fullAdder__1_2222 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2222

module PartialAdder__1_2223 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2129 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2132 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2135 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2138 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2141 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2144 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2147 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2150 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2153 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2156 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2159 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2162 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2165 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2168 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2171 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2174 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2177 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2180 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2183 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2186 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2189 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2192 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2195 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2198 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2201 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2204 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2207 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2210 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2213 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2216 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2219 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2222 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2223

module halfAdder__1_2032 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_2032

module fullAdder__1_2035 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2035

module fullAdder__1_2038 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2038

module fullAdder__1_2041 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2041

module fullAdder__1_2044 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_2044

module fullAdder__1_2047 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2047

module fullAdder__1_2050 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_2050

module fullAdder__1_2053 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_8), .A3 (n_0_4));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_4));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_2));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_8), .B2 (n_0_4));

endmodule //fullAdder__1_2053

module fullAdder__1_2056 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_2056

module fullAdder__1_2059 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (y));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (x), .A2 (n_0_5), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (sum), .A (n_0_0));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_2059

module fullAdder__1_2062 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2062

module fullAdder__1_2065 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


OAI21_X1 i_0_12 (.ZN (n_0_10), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (cout), .A1 (n_0_10), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_8), .A (y));
INV_X1 i_0_8 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_8), .A3 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_0 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_2065

module fullAdder__1_2068 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_2068

module fullAdder__1_2071 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2071

module fullAdder__1_2074 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2074

module fullAdder__1_2077 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2077

module fullAdder__1_2080 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2080

module fullAdder__1_2083 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2083

module fullAdder__1_2086 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2086

module fullAdder__1_2089 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2089

module fullAdder__1_2092 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2092

module fullAdder__1_2095 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2095

module fullAdder__1_2098 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2098

module fullAdder__1_2101 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2101

module fullAdder__1_2104 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2104

module fullAdder__1_2107 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2107

module fullAdder__1_2110 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2110

module fullAdder__1_2113 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2113

module fullAdder__1_2116 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2116

module fullAdder__1_2119 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2119

module fullAdder__1_2122 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2122

module fullAdder__1_2125 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2125

module PartialAdder__1_2126 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_2032 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_2035 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_2038 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_2041 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_2044 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_2047 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_2050 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_2053 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_2056 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_2059 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_2062 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_2065 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_2068 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_2071 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_2074 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_2077 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_2080 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_2083 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_2086 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_2089 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_2092 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_2095 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2098 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2101 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2104 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2107 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2110 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2113 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2116 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2119 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2122 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2125 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2126

module halfAdder__1_1935 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1935

module fullAdder__1_1938 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1938

module fullAdder__1_1941 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (n_0_4), .A3 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_3));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_5), .B1 (n_0_6), .B2 (n_0_3));

endmodule //fullAdder__1_1941

module fullAdder__1_1944 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1944

module fullAdder__1_1947 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1947

module fullAdder__1_1950 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1950

module fullAdder__1_1953 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;


OAI21_X1 i_0_4 (.ZN (n_0_2), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_1953

module fullAdder__1_1956 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1956

module fullAdder__1_1959 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_10), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (y), .A2 (cin));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_8), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1959

module fullAdder__1_1962 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1962

module fullAdder__1_1965 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1965

module fullAdder__1_1968 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1968

module fullAdder__1_1971 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1971

module fullAdder__1_1974 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1974

module fullAdder__1_1977 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1977

module fullAdder__1_1980 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1980

module fullAdder__1_1983 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1983

module fullAdder__1_1986 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1986

module fullAdder__1_1989 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1989

module fullAdder__1_1992 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1992

module fullAdder__1_1995 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1995

module fullAdder__1_1998 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1998

module fullAdder__1_2001 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2001

module fullAdder__1_2004 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2004

module fullAdder__1_2007 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2007

module fullAdder__1_2010 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2010

module fullAdder__1_2013 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2013

module fullAdder__1_2016 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2016

module fullAdder__1_2019 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2019

module fullAdder__1_2022 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2022

module fullAdder__1_2025 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2025

module fullAdder__1_2028 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_2028

module PartialAdder__1_2029 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1935 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1938 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1941 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1944 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1947 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1950 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1953 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1956 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1959 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1962 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1965 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1968 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1971 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1974 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1977 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1980 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1983 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1986 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1989 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1992 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1995 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1998 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_2001 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_2004 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_2007 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_2010 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_2013 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_2016 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_2019 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_2022 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_2025 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_2028 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_2029

module halfAdder__1_1838 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1838

module fullAdder__1_1841 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1841

module fullAdder__1_1844 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1844

module fullAdder__1_1847 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1847

module fullAdder__1_1850 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1850

module fullAdder__1_1853 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_0;
wire n_0_1;
wire n_0_2;


INV_X1 i_0_3 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NOR2_X1 i_0_8 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (x), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (x), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OR2_X1 i_0_4 (.ZN (n_0_3), .A1 (y), .A2 (cin));

endmodule //fullAdder__1_1853

module fullAdder__1_1856 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1856

module fullAdder__1_1859 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1859

module fullAdder__1_1862 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1862

module fullAdder__1_1865 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (sum), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_8 (.ZN (n_0_7), .A1 (n_0_3), .A2 (n_0_4), .A3 (n_0_1));
OAI21_X1 i_0_7 (.ZN (n_0_6), .A (y), .B1 (n_0_5), .B2 (n_0_2));
INV_X1 i_0_6 (.ZN (n_0_5), .A (n_0_1));
INV_X1 i_0_5 (.ZN (n_0_4), .A (y));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NOR2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_4));

endmodule //fullAdder__1_1865

module fullAdder__1_1868 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1868

module fullAdder__1_1871 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1871

module fullAdder__1_1874 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1874

module fullAdder__1_1877 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_5), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1877

module fullAdder__1_1880 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1880

module fullAdder__1_1883 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1883

module fullAdder__1_1886 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1886

module fullAdder__1_1889 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (cin));
NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (y), .A2 (n_0_11));
INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_9), .A2 (cin));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_10));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1889

module fullAdder__1_1892 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_7), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_7), .A3 (n_0_5));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1892

module fullAdder__1_1895 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1895

module fullAdder__1_1898 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1898

module fullAdder__1_1901 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1901

module fullAdder__1_1904 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1904

module fullAdder__1_1907 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1907

module fullAdder__1_1910 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1910

module fullAdder__1_1913 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1913

module fullAdder__1_1916 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1916

module fullAdder__1_1919 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1919

module fullAdder__1_1922 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1922

module fullAdder__1_1925 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1925

module fullAdder__1_1928 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1928

module fullAdder__1_1931 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1931

module PartialAdder__1_1932 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1838 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1841 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1844 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1847 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1850 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1853 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1856 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1859 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1862 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1865 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1868 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1871 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1874 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1877 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1880 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1883 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1886 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1889 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1892 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1895 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1898 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1901 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1904 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1907 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1910 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1913 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1916 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1919 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1922 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1925 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1928 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1931 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1932

module halfAdder__1_1741 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1741

module fullAdder__1_1744 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1744

module fullAdder__1_1747 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1747

module fullAdder__1_1750 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1750

module fullAdder__1_1753 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1753

module fullAdder__1_1756 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_1756

module fullAdder__1_1759 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (x));
INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_11), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1759

module fullAdder__1_1762 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_1762

module fullAdder__1_1765 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1765

module fullAdder__1_1768 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X2 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1768

module fullAdder__1_1771 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (x), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (x), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OR2_X1 i_0_4 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (x));
INV_X1 i_0_1 (.ZN (n_0_1), .A (cin));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_1771

module fullAdder__1_1774 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__1_1774

module fullAdder__1_1777 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_10), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (y), .A2 (cin));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_8), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_10));

endmodule //fullAdder__1_1777

module fullAdder__1_1780 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1780

module fullAdder__1_1783 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_8), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_3), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_5));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1783

module fullAdder__1_1786 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (y));
INV_X1 i_0_12 (.ZN (n_0_10), .A (x));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (n_0_10), .A2 (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_9), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_11), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_10), .A2 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_4));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));

endmodule //fullAdder__1_1786

module fullAdder__1_1789 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1789

module fullAdder__1_1792 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1792

module fullAdder__1_1795 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1795

module fullAdder__1_1798 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_10), .A3 (n_0_9));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1798

module fullAdder__1_1801 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1801

module fullAdder__1_1804 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1804

module fullAdder__1_1807 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1807

module fullAdder__1_1810 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1810

module fullAdder__1_1813 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1813

module fullAdder__1_1816 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1816

module fullAdder__1_1819 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1819

module fullAdder__1_1822 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1822

module fullAdder__1_1825 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1825

module fullAdder__1_1828 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1828

module fullAdder__1_1831 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1831

module fullAdder__1_1834 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1834

module PartialAdder__1_1835 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1741 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1744 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1747 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1750 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1753 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1756 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1759 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1762 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1765 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1768 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1771 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1774 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1777 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1780 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1783 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1786 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1789 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1792 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1795 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1798 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1801 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1804 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1807 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1810 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1813 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1816 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1819 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1822 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1825 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1828 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1831 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1834 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1835

module halfAdder__1_1644 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1644

module fullAdder__1_1647 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1647

module fullAdder__1_1650 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1650

module fullAdder__1_1653 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1653

module fullAdder__1_1656 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1656

module fullAdder__1_1659 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1659

module fullAdder__1_1662 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1662

module fullAdder__1_1665 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1665

module fullAdder__1_1668 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1668

module fullAdder__1_1671 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (y));
NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (n_0_11), .A2 (cin));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (y), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_10), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (x));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_11), .A2 (n_0_9));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_5), .A2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_6));
INV_X1 i_0_1 (.ZN (sum), .A (n_0_0));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_6), .A2 (n_0_4));

endmodule //fullAdder__1_1671

module fullAdder__1_1674 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


AOI21_X1 i_0_8 (.ZN (sum), .A (n_0_5), .B1 (y), .B2 (n_0_6));
OR2_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_3), .A2 (n_0_4));
NOR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_4), .A3 (y));
NOR2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1));
AND2_X1 i_0_3 (.ZN (n_0_3), .A1 (x), .A2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1674

module fullAdder__1_1677 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_5;
wire n_0_4;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_6;
wire n_0_7;
wire n_0_9;
wire n_0_8;
wire n_0_10;
wire n_0_11;
wire n_0_12;


INV_X1 i_0_14 (.ZN (n_0_12), .A (x));
INV_X1 i_0_13 (.ZN (n_0_11), .A (cin));
NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (y), .A2 (n_0_11));
INV_X1 i_0_11 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_9), .A1 (n_0_8), .A2 (cin));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_9), .A2 (n_0_10));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (n_0_12), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_2), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
INV_X1 i_0_4 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_3 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_5), .A1 (n_0_12), .A2 (n_0_11));
INV_X1 i_0_1 (.ZN (n_0_0), .A (n_0_5));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_4), .B1 (n_0_0), .B2 (n_0_8));

endmodule //fullAdder__1_1677

module fullAdder__1_1680 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1680

module fullAdder__1_1683 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1683

module fullAdder__1_1686 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1686

module fullAdder__1_1689 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_7), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_7), .A3 (n_0_5));
NAND2_X1 i_0_3 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_9), .B2 (n_0_0));

endmodule //fullAdder__1_1689

module fullAdder__1_1692 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


OAI21_X1 i_0_12 (.ZN (n_0_10), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (cout), .A1 (n_0_10), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_8), .A (y));
INV_X1 i_0_8 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_5), .A3 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_0 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_1692

module fullAdder__1_1695 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1695

module fullAdder__1_1698 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1698

module fullAdder__1_1701 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1701

module fullAdder__1_1704 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1704

module fullAdder__1_1707 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1707

module fullAdder__1_1710 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1710

module fullAdder__1_1713 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1713

module fullAdder__1_1716 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1716

module fullAdder__1_1719 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1719

module fullAdder__1_1722 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1722

module fullAdder__1_1725 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1725

module fullAdder__1_1728 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1728

module fullAdder__1_1731 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1731

module fullAdder__1_1734 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1734

module fullAdder__1_1737 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1737

module PartialAdder__1_1738 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1644 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1647 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1650 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1653 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1656 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1659 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1662 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1665 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1668 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1671 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1674 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1677 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1680 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1683 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1686 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1689 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1692 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1695 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1698 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1701 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1704 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1707 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1710 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1713 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1716 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1719 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1722 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1725 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1728 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1731 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1734 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1737 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1738

module halfAdder__1_1547 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1547

module fullAdder__1_1550 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1550

module fullAdder__1_1553 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1553

module fullAdder__1_1556 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1556

module fullAdder__1_1559 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1559

module fullAdder__1_1562 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1562

module fullAdder__1_1565 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1565

module fullAdder__1_1568 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1568

module fullAdder__1_1571 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1571

module fullAdder__1_1574 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1574

module fullAdder__1_1577 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1577

module fullAdder__1_1580 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


OAI21_X2 i_0_8 (.ZN (sum), .A (n_0_5), .B1 (n_0_6), .B2 (y));
AND2_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_3), .A2 (n_0_4));
NAND3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1));
OR2_X2 i_0_3 (.ZN (n_0_3), .A1 (x), .A2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1580

module fullAdder__1_1583 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_5), .B2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_4));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_1583

module fullAdder__1_1586 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1586

module fullAdder__1_1589 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1589

module fullAdder__1_1592 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1592

module fullAdder__1_1595 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1595

module fullAdder__1_1598 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1598

module fullAdder__1_1601 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (n_0_1));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_0), .A2 (cin));
NAND3_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (y), .A3 (n_0_9));
INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_0), .A2 (n_0_1));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_6), .A3 (n_0_5));
NAND2_X1 i_0_4 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_7));
NOR2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (cin));
OAI21_X1 i_0_2 (.ZN (cout), .A (n_0_5), .B1 (n_0_6), .B2 (n_0_2));
INV_X1 i_0_1 (.ZN (n_0_1), .A (cin));
INV_X1 i_0_0 (.ZN (n_0_0), .A (x));

endmodule //fullAdder__1_1601

module fullAdder__1_1604 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1604

module fullAdder__1_1607 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_1607

module fullAdder__1_1610 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (x));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9), .A3 (n_0_7));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_5));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1610

module fullAdder__1_1613 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1613

module fullAdder__1_1616 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1616

module fullAdder__1_1619 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1619

module fullAdder__1_1622 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1622

module fullAdder__1_1625 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1625

module fullAdder__1_1628 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1628

module fullAdder__1_1631 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1631

module fullAdder__1_1634 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1634

module fullAdder__1_1637 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1637

module fullAdder__1_1640 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1640

module PartialAdder__1_1641 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1547 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1550 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1553 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1556 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1559 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1562 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1565 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1568 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1571 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1574 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1577 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1580 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1583 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1586 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1589 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1592 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1595 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1598 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1601 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1604 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1607 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1610 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1613 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1616 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1619 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1622 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1625 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1628 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1631 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1634 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1637 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1640 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1641

module halfAdder__1_1450 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1450

module fullAdder__1_1453 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1453

module fullAdder__1_1456 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1456

module fullAdder__1_1459 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1459

module fullAdder__1_1462 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1462

module fullAdder__1_1465 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1465

module fullAdder__1_1468 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1468

module fullAdder__1_1471 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1471

module fullAdder__1_1474 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1474

module fullAdder__1_1477 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1477

module fullAdder__1_1480 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1480

module fullAdder__1_1483 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1483

module fullAdder__1_1486 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1486

module fullAdder__1_1489 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1489

module fullAdder__1_1492 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_0), .A2 (n_0_5));
AOI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (x), .B2 (cin));
OAI21_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3), .B1 (cin), .B2 (x));
OAI21_X1 i_0_3 (.ZN (sum), .A (n_0_2), .B1 (n_0_4), .B2 (n_0_6));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
INV_X1 i_0_1 (.ZN (n_0_0), .A (n_0_1));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_3), .A2 (n_0_5));

endmodule //fullAdder__1_1492

module fullAdder__1_1495 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_4), .B2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_2), .A (y));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_6));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1), .A3 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_6), .B1 (n_0_2), .B2 (n_0_5));

endmodule //fullAdder__1_1495

module fullAdder__1_1498 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1498

module fullAdder__1_1501 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_5), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1501

module fullAdder__1_1504 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1504

module fullAdder__1_1507 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1507

module fullAdder__1_1510 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
INV_X1 i_0_7 (.ZN (n_0_5), .A (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (y), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (x), .A3 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (x), .B1 (n_0_4), .B2 (n_0_3));
NOR2_X1 i_0_1 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_3));

endmodule //fullAdder__1_1510

module fullAdder__1_1513 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1513

module fullAdder__1_1516 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1516

module fullAdder__1_1519 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1519

module fullAdder__1_1522 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1522

module fullAdder__1_1525 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1525

module fullAdder__1_1528 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1528

module fullAdder__1_1531 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1531

module fullAdder__1_1534 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1534

module fullAdder__1_1537 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1537

module fullAdder__1_1540 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1540

module fullAdder__1_1543 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1543

module PartialAdder__1_1544 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1450 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1453 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1456 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1459 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1462 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1465 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1468 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1471 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1474 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1477 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1480 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1483 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1486 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1489 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1492 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1495 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1498 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1501 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1504 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1507 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1510 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1513 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1516 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1519 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1522 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1525 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1528 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1531 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1534 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1537 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1540 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1543 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1544

module halfAdder__1_1353 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1353

module fullAdder__1_1356 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1356

module fullAdder__1_1359 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1359

module fullAdder__1_1362 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1362

module fullAdder__1_1365 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1365

module fullAdder__1_1368 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1368

module fullAdder__1_1371 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1371

module fullAdder__1_1374 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1374

module fullAdder__1_1377 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1377

module fullAdder__1_1380 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1380

module fullAdder__1_1383 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1383

module fullAdder__1_1386 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1386

module fullAdder__1_1389 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1389

module fullAdder__1_1392 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1392

module fullAdder__1_1395 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_10), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (y), .A2 (cin));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_8), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1395

module fullAdder__1_1398 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (y), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (y));
INV_X1 i_0_5 (.ZN (n_0_3), .A (cin));
INV_X1 i_0_4 (.ZN (n_0_2), .A (x));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_3));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_4), .A3 (n_0_8));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_6), .B1 (n_0_4), .B2 (n_0_8));

endmodule //fullAdder__1_1398

module fullAdder__1_1401 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (n_0_8));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_7), .A3 (n_0_5));
NAND2_X1 i_0_3 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_9), .B2 (n_0_0));

endmodule //fullAdder__1_1401

module fullAdder__1_1404 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1404

module fullAdder__1_1407 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1407

module fullAdder__1_1410 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1410

module fullAdder__1_1413 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1413

module fullAdder__1_1416 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1416

module fullAdder__1_1419 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1419

module fullAdder__1_1422 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
NOR2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_10), .A2 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_8));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1422

module fullAdder__1_1425 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1425

module fullAdder__1_1428 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1428

module fullAdder__1_1431 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1431

module fullAdder__1_1434 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1434

module fullAdder__1_1437 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1437

module fullAdder__1_1440 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1440

module fullAdder__1_1443 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1443

module fullAdder__1_1446 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1446

module PartialAdder__1_1447 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1353 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1356 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1359 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1362 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1365 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1368 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1371 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1374 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1377 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1380 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1383 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1386 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1389 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1392 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1395 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1398 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1401 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1404 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1407 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1410 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1413 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1416 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1419 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1422 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1425 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1428 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1431 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1434 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1437 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1440 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1443 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1446 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1447

module halfAdder__1_1256 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1256

module fullAdder__1_1259 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1259

module fullAdder__1_1262 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1262

module fullAdder__1_1265 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1265

module fullAdder__1_1268 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1268

module fullAdder__1_1271 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1271

module fullAdder__1_1274 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1274

module fullAdder__1_1277 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1277

module fullAdder__1_1280 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1280

module fullAdder__1_1283 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1283

module fullAdder__1_1286 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1286

module fullAdder__1_1289 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1289

module fullAdder__1_1292 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (x), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (x), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OR2_X1 i_0_4 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (x));
INV_X1 i_0_1 (.ZN (n_0_1), .A (cin));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_1292

module fullAdder__1_1295 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_6 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (x), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (x), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (cin));
OR2_X2 i_0_0 (.ZN (n_0_0), .A1 (y), .A2 (cin));

endmodule //fullAdder__1_1295

module fullAdder__1_1298 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X2 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1298

module fullAdder__1_1301 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (n_0_1));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_1));
NAND2_X1 i_0_8 (.ZN (sum), .A1 (n_0_7), .A2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (y), .A2 (n_0_6));
INV_X1 i_0_5 (.ZN (n_0_4), .A (y));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (n_0_4), .A2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1301

module fullAdder__1_1304 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


INV_X1 i_0_13 (.ZN (n_0_11), .A (x));
NOR2_X1 i_0_12 (.ZN (n_0_10), .A1 (y), .A2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (n_0_9));
OAI21_X1 i_0_9 (.ZN (n_0_7), .A (n_0_11), .B1 (n_0_8), .B2 (n_0_10));
INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
INV_X1 i_0_7 (.ZN (n_0_5), .A (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (x), .A3 (n_0_9));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_1304

module fullAdder__1_1307 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1307

module fullAdder__1_1310 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1310

module fullAdder__1_1313 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_1313

module fullAdder__1_1316 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1316

module fullAdder__1_1319 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1319

module fullAdder__1_1322 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


AOI21_X1 i_0_9 (.ZN (sum), .A (n_0_6), .B1 (n_0_7), .B2 (x));
OR2_X1 i_0_8 (.ZN (n_0_7), .A1 (n_0_4), .A2 (n_0_5));
NOR3_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_4), .A2 (n_0_5), .A3 (x));
NOR2_X1 i_0_6 (.ZN (n_0_5), .A1 (y), .A2 (n_0_3));
AND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (n_0_3));
INV_X1 i_0_4 (.ZN (n_0_3), .A (cin));
INV_X1 i_0_3 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));

endmodule //fullAdder__1_1322

module fullAdder__1_1325 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1325

module fullAdder__1_1328 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1328

module fullAdder__1_1331 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (n_0_4), .A3 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_3));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_5), .B1 (n_0_6), .B2 (n_0_3));

endmodule //fullAdder__1_1331

module fullAdder__1_1334 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1334

module fullAdder__1_1337 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1337

module fullAdder__1_1340 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1340

module fullAdder__1_1343 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1343

module fullAdder__1_1346 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1346

module fullAdder__1_1349 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1349

module PartialAdder__1_1350 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1256 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1259 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1262 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1265 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1268 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1271 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1274 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1277 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1280 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1283 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1286 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1289 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1292 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1295 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1298 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1301 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1304 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1307 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1310 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1313 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1316 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1319 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1322 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1325 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1328 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1331 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1334 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1337 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1340 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1343 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1346 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1349 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1350

module halfAdder__1_1159 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1159

module fullAdder__1_1162 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1162

module fullAdder__1_1165 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1165

module fullAdder__1_1168 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1168

module fullAdder__1_1171 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1171

module fullAdder__1_1174 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1174

module fullAdder__1_1177 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1177

module fullAdder__1_1180 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1180

module fullAdder__1_1183 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1183

module fullAdder__1_1186 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1186

module fullAdder__1_1189 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1189

module fullAdder__1_1192 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1192

module fullAdder__1_1195 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X2 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__1_1195

module fullAdder__1_1198 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1198

module fullAdder__1_1201 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1201

module fullAdder__1_1204 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (x));
INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (y), .A2 (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_10), .A2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7), .A3 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_1204

module fullAdder__1_1207 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1207

module fullAdder__1_1210 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1210

module fullAdder__1_1213 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1213

module fullAdder__1_1216 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1216

module fullAdder__1_1219 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1219

module fullAdder__1_1222 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1222

module fullAdder__1_1225 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1225

module fullAdder__1_1228 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1228

module fullAdder__1_1231 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1231

module fullAdder__1_1234 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_10), .A2 (n_0_7), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1234

module fullAdder__1_1237 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1237

module fullAdder__1_1240 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1240

module fullAdder__1_1243 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1243

module fullAdder__1_1246 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1246

module fullAdder__1_1249 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1249

module fullAdder__1_1252 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1252

module PartialAdder__1_1253 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1159 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1162 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1165 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1168 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1171 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1174 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1177 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1180 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1183 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1186 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1189 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1192 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1195 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1198 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1201 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1204 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1207 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1210 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1213 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1216 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1219 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1222 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1225 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1228 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1231 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1234 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1237 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1240 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1243 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1246 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1249 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1252 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1253

module halfAdder__1_1062 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_1062

module fullAdder__1_1065 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1065

module fullAdder__1_1068 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1068

module fullAdder__1_1071 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1071

module fullAdder__1_1074 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1074

module fullAdder__1_1077 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1077

module fullAdder__1_1080 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1080

module fullAdder__1_1083 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1083

module fullAdder__1_1086 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1086

module fullAdder__1_1089 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1089

module fullAdder__1_1092 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1092

module fullAdder__1_1095 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1095

module fullAdder__1_1098 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1098

module fullAdder__1_1101 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X2 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1101

module fullAdder__1_1104 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1104

module fullAdder__1_1107 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X2 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_1107

module fullAdder__1_1110 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_6));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_5), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_1110

module fullAdder__1_1113 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_0), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
AOI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (y));
NOR2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_1113

module fullAdder__1_1116 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_1116

module fullAdder__1_1119 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


OAI21_X1 i_0_12 (.ZN (n_0_10), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (cout), .A1 (n_0_10), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_8), .A (y));
INV_X1 i_0_8 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_5), .A3 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y), .A3 (n_0_2));
NAND2_X2 i_0_0 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_1119

module fullAdder__1_1122 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1122

module fullAdder__1_1125 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1125

module fullAdder__1_1128 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1128

module fullAdder__1_1131 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1131

module fullAdder__1_1134 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1134

module fullAdder__1_1137 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1137

module fullAdder__1_1140 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NOR2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (n_0_10));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (n_0_10));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
OAI21_X1 i_0_8 (.ZN (n_0_6), .A (y), .B1 (n_0_7), .B2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_5), .A (y));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_4));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
OAI21_X1 i_0_3 (.ZN (n_0_1), .A (n_0_5), .B1 (n_0_3), .B2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_6), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (sum), .A (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_5), .B2 (n_0_4));

endmodule //fullAdder__1_1140

module fullAdder__1_1143 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1143

module fullAdder__1_1146 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1146

module fullAdder__1_1149 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1149

module fullAdder__1_1152 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1152

module fullAdder__1_1155 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1155

module PartialAdder__1_1156 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_1062 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_1065 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_1068 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_1071 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_1074 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_1077 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_1080 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_1083 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_1086 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_1089 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_1092 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_1095 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1098 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1101 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1104 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1107 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1110 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1113 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1116 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1119 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1122 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1125 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1128 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1131 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1134 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1137 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1140 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1143 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1146 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1149 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1152 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1155 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1156

module halfAdder__1_965 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_965

module fullAdder__1_968 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_968

module fullAdder__1_971 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_971

module fullAdder__1_974 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_974

module fullAdder__1_977 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_977

module fullAdder__1_980 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_980

module fullAdder__1_983 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_983

module fullAdder__1_986 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_986

module fullAdder__1_989 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_989

module fullAdder__1_992 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_992

module fullAdder__1_995 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_995

module fullAdder__1_998 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_998

module fullAdder__1_1001 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1001

module fullAdder__1_1004 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1004

module fullAdder__1_1007 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_0;
wire n_0_1;
wire n_0_3;
wire n_0_5;
wire n_0_2;
wire n_0_9;
wire n_0_4;


NAND2_X1 i_0_11 (.ZN (n_0_4), .A1 (x), .A2 (cin));
INV_X1 i_0_10 (.ZN (n_0_9), .A (n_0_4));
NOR2_X1 i_0_7 (.ZN (n_0_2), .A1 (x), .A2 (cin));
OAI21_X1 i_0_6 (.ZN (n_0_5), .A (y), .B1 (n_0_9), .B2 (n_0_2));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (n_0_7));
AOI21_X1 i_0_4 (.ZN (n_0_1), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_3 (.ZN (n_0_0), .A1 (n_0_3), .A2 (n_0_1));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_0));
INV_X1 i_0_1 (.ZN (n_0_8), .A (y));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_8), .B2 (n_0_4));

endmodule //fullAdder__1_1007

module fullAdder__1_1010 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1010

module fullAdder__1_1013 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1013

module fullAdder__1_1016 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1016

module fullAdder__1_1019 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NOR2_X2 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_5), .B2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_4));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_1019

module fullAdder__1_1022 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_5), .B2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_4));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_1022

module fullAdder__1_1025 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (n_0_9));
NOR2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (n_0_10));
OAI21_X1 i_0_8 (.ZN (n_0_6), .A (y), .B1 (n_0_8), .B2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (y));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_4));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
OAI21_X1 i_0_3 (.ZN (n_0_1), .A (n_0_5), .B1 (n_0_3), .B2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_6), .A2 (n_0_1));
INV_X2 i_0_1 (.ZN (sum), .A (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_5), .B2 (n_0_4));

endmodule //fullAdder__1_1025

module fullAdder__1_1028 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1028

module fullAdder__1_1031 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1031

module fullAdder__1_1034 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_1034

module fullAdder__1_1037 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1037

module fullAdder__1_1040 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (y));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (x), .A2 (n_0_5), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (sum), .A (n_0_0));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_1), .A2 (n_0_4));

endmodule //fullAdder__1_1040

module fullAdder__1_1043 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1043

module fullAdder__1_1046 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1046

module fullAdder__1_1049 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1049

module fullAdder__1_1052 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1052

module fullAdder__1_1055 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1055

module fullAdder__1_1058 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_1058

module PartialAdder__1_1059 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_965 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_968 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_971 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_974 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_977 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_980 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_983 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_986 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_989 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_992 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_995 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_998 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_1001 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_1004 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_1007 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_1010 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_1013 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_1016 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_1019 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_1022 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_1025 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_1028 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_1031 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_1034 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_1037 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_1040 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_1043 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_1046 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_1049 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_1052 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_1055 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_1058 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_1059

module halfAdder__1_868 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_868

module fullAdder__1_871 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_871

module fullAdder__1_874 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_874

module fullAdder__1_877 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_877

module fullAdder__1_880 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_880

module fullAdder__1_883 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_883

module fullAdder__1_886 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_886

module fullAdder__1_889 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_889

module fullAdder__1_892 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_892

module fullAdder__1_895 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_895

module fullAdder__1_898 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_898

module fullAdder__1_901 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_901

module fullAdder__1_904 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_904

module fullAdder__1_907 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_907

module fullAdder__1_910 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_910

module fullAdder__1_913 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_913

module fullAdder__1_916 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_6 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (x), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (x), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (cin));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (y), .A2 (cin));

endmodule //fullAdder__1_916

module fullAdder__1_919 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_919

module fullAdder__1_922 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__1_922

module fullAdder__1_925 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X2 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_925

module fullAdder__1_928 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_7;
wire n_0_8;


AOI22_X1 i_0_10 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_8), .B1 (x), .B2 (n_0_7));
INV_X1 i_0_9 (.ZN (n_0_8), .A (n_0_7));
NAND2_X1 i_0_8 (.ZN (n_0_7), .A1 (n_0_1), .A2 (n_0_0));
OAI21_X1 i_0_7 (.ZN (cout), .A (n_0_4), .B1 (n_0_5), .B2 (n_0_2));
INV_X1 i_0_5 (.ZN (n_0_5), .A (x));
OAI21_X1 i_0_4 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
INV_X1 i_0_3 (.ZN (n_0_3), .A (y));
INV_X1 i_0_2 (.ZN (n_0_2), .A (cin));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (n_0_2));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (n_0_3), .A2 (cin));

endmodule //fullAdder__1_928

module fullAdder__1_931 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_931

module fullAdder__1_934 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_934

module fullAdder__1_937 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_937

module fullAdder__1_940 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_8), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_940

module fullAdder__1_943 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_943

module fullAdder__1_946 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


NOR2_X1 i_0_12 (.ZN (n_0_10), .A1 (x), .A2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
OAI21_X1 i_0_10 (.ZN (cout), .A (n_0_9), .B1 (n_0_10), .B2 (n_0_8));
INV_X1 i_0_9 (.ZN (n_0_8), .A (y));
INV_X1 i_0_8 (.ZN (n_0_7), .A (cin));
NOR2_X1 i_0_7 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_5));
OAI21_X1 i_0_4 (.ZN (n_0_3), .A (n_0_8), .B1 (n_0_4), .B2 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_2), .A (x));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_2), .A2 (cin));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y), .A3 (n_0_5));
NAND2_X1 i_0_0 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_946

module fullAdder__1_949 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_949

module fullAdder__1_952 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_952

module fullAdder__1_955 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_955

module fullAdder__1_958 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_958

module fullAdder__1_961 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_961

module PartialAdder__1_962 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_868 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_871 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_874 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_877 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_880 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_883 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_886 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_889 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_892 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_895 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_898 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_901 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_904 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_907 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_910 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_913 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_916 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_919 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_922 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_925 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_928 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_931 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_934 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_937 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_940 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_943 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_946 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_949 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_952 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_955 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_958 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_961 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_962

module halfAdder__1_771 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_771

module fullAdder__1_774 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_774

module fullAdder__1_777 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_777

module fullAdder__1_780 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_780

module fullAdder__1_783 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_783

module fullAdder__1_786 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_786

module fullAdder__1_789 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_789

module fullAdder__1_792 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_792

module fullAdder__1_795 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_795

module fullAdder__1_798 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_798

module fullAdder__1_801 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_801

module fullAdder__1_804 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_804

module fullAdder__1_807 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_807

module fullAdder__1_810 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_810

module fullAdder__1_813 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_813

module fullAdder__1_816 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_816

module fullAdder__1_819 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_819

module fullAdder__1_822 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_822

module fullAdder__1_825 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X2 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_825

module fullAdder__1_828 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NOR2_X1 i_0_9 (.ZN (sum), .A1 (n_0_6), .A2 (n_0_7));
AOI21_X1 i_0_8 (.ZN (n_0_7), .A (x), .B1 (n_0_5), .B2 (n_0_4));
AND3_X1 i_0_7 (.ZN (n_0_6), .A1 (n_0_4), .A2 (x), .A3 (n_0_5));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (y), .A2 (cin));
OR2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (cin));
OR2_X1 i_0_4 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (n_0_3), .B1 (n_0_1), .B2 (y));
INV_X1 i_0_0 (.ZN (cout), .A (n_0_0));

endmodule //fullAdder__1_828

module fullAdder__1_831 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_831

module fullAdder__1_834 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__1_834

module fullAdder__1_837 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_837

module fullAdder__1_840 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_840

module fullAdder__1_843 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_843

module fullAdder__1_846 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_8), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_3), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_5));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_846

module fullAdder__1_849 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_849

module fullAdder__1_852 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


OAI21_X1 i_0_12 (.ZN (n_0_10), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (x), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (cout), .A1 (n_0_10), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_8), .A (y));
INV_X1 i_0_8 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_5), .A3 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_0 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_852

module fullAdder__1_855 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_855

module fullAdder__1_858 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_858

module fullAdder__1_861 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_861

module fullAdder__1_864 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_864

module PartialAdder__1_865 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_771 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_774 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_777 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_780 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_783 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_786 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_789 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_792 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_795 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_798 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_801 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_804 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_807 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_810 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_813 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_816 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_819 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_822 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_825 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_828 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_831 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_834 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_837 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_840 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_843 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_846 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_849 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_852 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_855 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_858 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_861 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_864 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_865

module halfAdder__1_674 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_674

module fullAdder__1_677 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_677

module fullAdder__1_680 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_680

module fullAdder__1_683 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_683

module fullAdder__1_686 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_686

module fullAdder__1_689 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_689

module fullAdder__1_692 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_692

module fullAdder__1_695 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_695

module fullAdder__1_698 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_698

module fullAdder__1_701 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_701

module fullAdder__1_704 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_704

module fullAdder__1_707 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_707

module fullAdder__1_710 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_710

module fullAdder__1_713 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_713

module fullAdder__1_716 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_716

module fullAdder__1_719 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_719

module fullAdder__1_722 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_722

module fullAdder__1_725 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_725

module fullAdder__1_728 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_728

module fullAdder__1_731 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


AOI22_X1 i_0_8 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_6), .B1 (x), .B2 (n_0_5));
INV_X1 i_0_7 (.ZN (n_0_6), .A (n_0_5));
OAI22_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (cin), .B1 (y), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (cin));
INV_X1 i_0_3 (.ZN (n_0_3), .A (y));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_731

module fullAdder__1_734 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
XNOR2_X1 i_0_7 (.ZN (n_0_5), .A (y), .B (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_734

module fullAdder__1_737 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


AOI22_X1 i_0_10 (.ZN (sum), .A1 (n_0_6), .A2 (n_0_8), .B1 (x), .B2 (n_0_7));
INV_X1 i_0_9 (.ZN (n_0_8), .A (n_0_7));
NAND2_X1 i_0_8 (.ZN (n_0_7), .A1 (n_0_1), .A2 (n_0_4));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
INV_X1 i_0_6 (.ZN (n_0_5), .A (cin));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (n_0_5));
INV_X1 i_0_3 (.ZN (n_0_3), .A (y));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_3), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_737

module fullAdder__1_740 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_740

module fullAdder__1_743 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_743

module fullAdder__1_746 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_746

module fullAdder__1_749 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_8), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_3), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_5));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_749

module fullAdder__1_752 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_5), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_752

module fullAdder__1_755 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (n_0_4), .A3 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_3));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_0));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_5), .B1 (n_0_6), .B2 (n_0_3));

endmodule //fullAdder__1_755

module fullAdder__1_758 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


INV_X1 i_0_7 (.ZN (n_0_5), .A (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (x));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_758

module fullAdder__1_761 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_761

module fullAdder__1_764 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_764

module fullAdder__1_767 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_767

module PartialAdder__1_768 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_674 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_677 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_680 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_683 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_686 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_689 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_692 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_695 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_698 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_701 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_704 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_707 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_710 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_713 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_716 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_719 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_722 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_725 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_728 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_731 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_734 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_737 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_740 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_743 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_746 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_749 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_752 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_755 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_758 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_761 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_764 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_767 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_768

module halfAdder__1_577 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_577

module fullAdder__1_580 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_580

module fullAdder__1_583 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_583

module fullAdder__1_586 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_586

module fullAdder__1_589 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_589

module fullAdder__1_592 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_592

module fullAdder__1_595 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_595

module fullAdder__1_598 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_598

module fullAdder__1_601 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_601

module fullAdder__1_604 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_604

module fullAdder__1_607 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_607

module fullAdder__1_610 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_610

module fullAdder__1_613 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_613

module fullAdder__1_616 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_616

module fullAdder__1_619 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_619

module fullAdder__1_622 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_622

module fullAdder__1_625 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_625

module fullAdder__1_628 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_0), .A2 (n_0_5));
AOI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (x), .B2 (cin));
OAI21_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3), .B1 (cin), .B2 (x));
OAI21_X1 i_0_3 (.ZN (sum), .A (n_0_2), .B1 (n_0_4), .B2 (n_0_6));
NOR2_X1 i_0_2 (.ZN (cout), .A1 (n_0_3), .A2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
INV_X1 i_0_0 (.ZN (n_0_0), .A (n_0_1));

endmodule //fullAdder__1_628

module fullAdder__1_631 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_631

module fullAdder__1_634 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_634

module fullAdder__1_637 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_637

module fullAdder__1_640 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_640

module fullAdder__1_643 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (y), .B1 (n_0_7), .B2 (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_0), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));
INV_X1 i_0_1 (.ZN (n_0_1), .A (cin));
INV_X1 i_0_0 (.ZN (n_0_0), .A (x));

endmodule //fullAdder__1_643

module fullAdder__1_646 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (y), .B1 (x), .B2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y), .B1 (n_0_1), .B2 (n_0_6));
NAND2_X2 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_4), .A2 (n_0_6));

endmodule //fullAdder__1_646

module fullAdder__1_649 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_649

module fullAdder__1_652 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_652

module fullAdder__1_655 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_6), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_655

module fullAdder__1_658 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_658

module fullAdder__1_661 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_6));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_7), .A3 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_7));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_4));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_7));

endmodule //fullAdder__1_661

module fullAdder__1_664 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


OR2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_664

module fullAdder__1_667 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_667

module fullAdder__1_670 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_670

module PartialAdder__1_671 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_577 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_580 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_583 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_586 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_589 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_592 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_595 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_598 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_601 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_604 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_607 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_610 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_613 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_616 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_619 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_622 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_625 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_628 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_631 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_634 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_637 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_640 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_643 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_646 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_649 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_652 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_655 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_658 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_661 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_664 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_667 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_670 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_671

module halfAdder__1_480 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_480

module fullAdder__1_483 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_483

module fullAdder__1_486 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_486

module fullAdder__1_489 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_489

module fullAdder__1_492 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_492

module fullAdder__1_495 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_495

module fullAdder__1_498 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_498

module fullAdder__1_501 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_501

module fullAdder__1_504 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_504

module fullAdder__1_507 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_507

module fullAdder__1_510 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_510

module fullAdder__1_513 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_513

module fullAdder__1_516 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_516

module fullAdder__1_519 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_519

module fullAdder__1_522 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_522

module fullAdder__1_525 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_525

module fullAdder__1_528 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_528

module fullAdder__1_531 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_531

module fullAdder__1_534 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_534

module fullAdder__1_537 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


OAI21_X1 i_0_7 (.ZN (n_0_5), .A (n_0_0), .B1 (cin), .B2 (x));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
OAI21_X1 i_0_3 (.ZN (n_0_1), .A (y), .B1 (n_0_2), .B2 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_5));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_4));

endmodule //fullAdder__1_537

module fullAdder__1_540 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_540

module fullAdder__1_543 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X2 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_543

module fullAdder__1_546 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_546

module fullAdder__1_549 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_6));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_5), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_549

module fullAdder__1_552 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_552

module fullAdder__1_555 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_555

module fullAdder__1_558 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_558

module fullAdder__1_561 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (n_0_9));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_561

module fullAdder__1_564 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NOR2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (n_0_9));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (n_0_10), .B1 (n_0_6), .B2 (n_0_8));
INV_X1 i_0_6 (.ZN (n_0_4), .A (x));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_7));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_564

module fullAdder__1_567 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (y), .B1 (n_0_4), .B2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_2), .A (y));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_6));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1), .A3 (n_0_5));
NAND2_X1 i_0_1 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_3));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_6), .B1 (n_0_2), .B2 (n_0_5));

endmodule //fullAdder__1_567

module fullAdder__1_570 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


OR2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_570

module fullAdder__1_573 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_573

module PartialAdder__1_574 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_480 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_483 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_486 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_489 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_492 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_495 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_498 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_501 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_504 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_507 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_510 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_513 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_516 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_519 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_522 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_525 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_528 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_531 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_534 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_537 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_540 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_543 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_546 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_549 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_552 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_555 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_558 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_561 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_564 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_567 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_570 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_573 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_574

module halfAdder__1_383 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_383

module fullAdder__1_386 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_386

module fullAdder__1_389 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_389

module fullAdder__1_392 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_392

module fullAdder__1_395 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_395

module fullAdder__1_398 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_398

module fullAdder__1_401 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_401

module fullAdder__1_404 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_404

module fullAdder__1_407 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_407

module fullAdder__1_410 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_410

module fullAdder__1_413 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_413

module fullAdder__1_416 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_416

module fullAdder__1_419 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_419

module fullAdder__1_422 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_422

module fullAdder__1_425 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_425

module fullAdder__1_428 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_428

module fullAdder__1_431 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_431

module fullAdder__1_434 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_434

module fullAdder__1_437 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_3), .B2 (n_0_1));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_437

module fullAdder__1_440 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_440

module fullAdder__1_443 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_443

module fullAdder__1_446 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_446

module fullAdder__1_449 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_449

module fullAdder__1_452 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (x), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (x), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (cin));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (y), .A2 (cin));

endmodule //fullAdder__1_452

module fullAdder__1_455 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
XNOR2_X1 i_0_7 (.ZN (n_0_5), .A (y), .B (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_455

module fullAdder__1_458 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_458

module fullAdder__1_461 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_461

module fullAdder__1_464 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_464

module fullAdder__1_467 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (n_0_6), .A2 (n_0_4));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (n_0_10));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
NAND2_X1 i_0_9 (.ZN (cout), .A1 (n_0_9), .A2 (n_0_8));
INV_X1 i_0_8 (.ZN (n_0_7), .A (y));
INV_X1 i_0_7 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_6), .A2 (cin));
INV_X1 i_0_5 (.ZN (n_0_4), .A (cin));
NAND2_X1 i_0_4 (.ZN (n_0_3), .A1 (x), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (n_0_5), .A2 (n_0_3));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_7));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_5), .A3 (n_0_3));
NAND2_X1 i_0_0 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_0));

endmodule //fullAdder__1_467

module fullAdder__1_470 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_5), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_470

module fullAdder__1_473 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_473

module fullAdder__1_476 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


OR2_X1 i_0_5 (.ZN (n_0_3), .A1 (cin), .A2 (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (y), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (cin), .A2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_476

module PartialAdder__1_477 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_383 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_386 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_389 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_392 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_395 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_398 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_401 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_404 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_407 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_410 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_413 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_416 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_419 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_422 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_425 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_428 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_431 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_434 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_437 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_440 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_443 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_446 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_449 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_452 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_455 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_458 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_461 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_464 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_467 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_470 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_473 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_476 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_477

module halfAdder__1_286 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_286

module fullAdder__1_289 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_289

module fullAdder__1_292 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_292

module fullAdder__1_295 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_295

module fullAdder__1_298 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_298

module fullAdder__1_301 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_301

module fullAdder__1_304 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_304

module fullAdder__1_307 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_307

module fullAdder__1_310 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_310

module fullAdder__1_313 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_313

module fullAdder__1_316 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_316

module fullAdder__1_319 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_319

module fullAdder__1_322 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_322

module fullAdder__1_325 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_325

module fullAdder__1_328 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_328

module fullAdder__1_331 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_331

module fullAdder__1_334 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_334

module fullAdder__1_337 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_337

module fullAdder__1_340 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_340

module fullAdder__1_343 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_343

module fullAdder__1_346 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (y));
INV_X1 i_0_8 (.ZN (n_0_6), .A (cin));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (y), .A2 (cin));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (x), .A3 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (x), .B1 (n_0_5), .B2 (n_0_4));
NOR2_X1 i_0_2 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_3), .A2 (n_0_0));

endmodule //fullAdder__1_346

module fullAdder__1_349 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_4 (.ZN (n_0_3), .A (y), .B (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (x));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_349

module fullAdder__1_352 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_352

module fullAdder__1_355 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (y));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (cin));
OAI21_X1 i_0_5 (.ZN (cout), .A (n_0_4), .B1 (n_0_5), .B2 (n_0_6));
NOR2_X2 i_0_4 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_3));
AOI21_X1 i_0_3 (.ZN (n_0_3), .A (x), .B1 (n_0_0), .B2 (n_0_1));
AND3_X1 i_0_2 (.ZN (n_0_2), .A1 (x), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (cin));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (y), .A2 (cin));

endmodule //fullAdder__1_355

module fullAdder__1_358 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


AOI22_X1 i_0_8 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_5), .B1 (x), .B2 (n_0_6));
INV_X1 i_0_7 (.ZN (n_0_6), .A (n_0_5));
NAND2_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_4), .A2 (n_0_1));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
OAI21_X1 i_0_4 (.ZN (cout), .A (n_0_1), .B1 (n_0_0), .B2 (n_0_3));
NOR2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (y), .A2 (cin));
INV_X1 i_0_0 (.ZN (n_0_0), .A (x));

endmodule //fullAdder__1_358

module fullAdder__1_361 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (x));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_6));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_361

module fullAdder__1_364 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (y));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (y), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (x), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_4));
AOI21_X1 i_0_4 (.ZN (n_0_2), .A (x), .B1 (n_0_6), .B2 (n_0_5));
NOR2_X1 i_0_3 (.ZN (sum), .A1 (n_0_3), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_7), .B2 (n_0_1));

endmodule //fullAdder__1_364

module fullAdder__1_367 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_9), .A2 (n_0_6), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_8));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_367

module fullAdder__1_370 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_370

module fullAdder__1_373 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_373

module fullAdder__1_376 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_9), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (y), .A2 (n_0_4));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (n_0_6));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_376

module fullAdder__1_379 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_379

module PartialAdder__1_380 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_286 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_289 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_292 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_295 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_298 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_301 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_304 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_307 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_310 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_313 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_316 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_319 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_322 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_325 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_328 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_331 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_334 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_337 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_340 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_343 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_346 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_349 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_352 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_355 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_358 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_361 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_364 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_367 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_370 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_373 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_376 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_379 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_380

module halfAdder__1_189 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_189

module fullAdder__1_192 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_192

module fullAdder__1_195 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_195

module fullAdder__1_198 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_198

module fullAdder__1_201 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_201

module fullAdder__1_204 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_204

module fullAdder__1_207 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_207

module fullAdder__1_210 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_210

module fullAdder__1_213 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_213

module fullAdder__1_216 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_216

module fullAdder__1_219 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_219

module fullAdder__1_222 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_222

module fullAdder__1_225 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_225

module fullAdder__1_228 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_228

module fullAdder__1_231 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_231

module fullAdder__1_234 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_234

module fullAdder__1_237 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_237

module fullAdder__1_240 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_240

module fullAdder__1_243 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (y));
INV_X1 i_0_11 (.ZN (n_0_9), .A (cin));
NOR2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (x), .A2 (n_0_9));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (n_0_10), .B1 (n_0_6), .B2 (n_0_8));
INV_X1 i_0_6 (.ZN (n_0_4), .A (x));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_7));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_243

module fullAdder__1_246 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_246

module fullAdder__1_249 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_249

module fullAdder__1_252 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_11;
wire n_0_12;


NOR2_X1 i_0_14 (.ZN (n_0_12), .A1 (y), .A2 (cin));
NAND2_X1 i_0_13 (.ZN (n_0_11), .A1 (n_0_0), .A2 (n_0_12));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (cin));
INV_X1 i_0_10 (.ZN (n_0_8), .A (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_0), .A2 (n_0_8));
OR2_X1 i_0_8 (.ZN (n_0_6), .A1 (y), .A2 (cin));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (n_0_9), .A3 (n_0_6));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_11), .A2 (n_0_7), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (sum), .A (n_0_4));
NOR2_X1 i_0_4 (.ZN (n_0_3), .A1 (x), .A2 (cin));
AOI21_X1 i_0_3 (.ZN (n_0_2), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_2 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_3));
INV_X1 i_0_0 (.ZN (n_0_0), .A (x));

endmodule //fullAdder__1_252

module fullAdder__1_255 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_4 (.ZN (n_0_3), .A (y), .B (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (x));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_255

module fullAdder__1_258 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_258

module fullAdder__1_261 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X2 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_261

module fullAdder__1_264 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (sum), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
NOR2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_1));

endmodule //fullAdder__1_264

module fullAdder__1_267 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_267

module fullAdder__1_270 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (x));
NOR2_X1 i_0_11 (.ZN (n_0_9), .A1 (y), .A2 (cin));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (y), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (n_0_8));
OAI21_X1 i_0_8 (.ZN (n_0_6), .A (n_0_10), .B1 (n_0_7), .B2 (n_0_9));
INV_X1 i_0_7 (.ZN (n_0_5), .A (y));
INV_X1 i_0_6 (.ZN (n_0_4), .A (cin));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (x), .A3 (n_0_8));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_4), .B2 (n_0_10));

endmodule //fullAdder__1_270

module fullAdder__1_273 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (x), .A2 (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (n_0_7));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_9), .A3 (n_0_8));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (cin));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (y), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_5), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_8));

endmodule //fullAdder__1_273

module fullAdder__1_276 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_1), .A2 (x), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_276

module fullAdder__1_279 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (y));
INV_X1 i_0_10 (.ZN (n_0_8), .A (cin));
INV_X1 i_0_9 (.ZN (n_0_7), .A (x));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (x), .A2 (cin));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_9), .A3 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_8));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (y), .A3 (n_0_2));
NAND2_X1 i_0_2 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_6), .A2 (y));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_5));

endmodule //fullAdder__1_279

module fullAdder__1_282 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OAI21_X1 i_0_6 (.ZN (n_0_5), .A (y), .B1 (n_0_1), .B2 (n_0_3));
OR3_X1 i_0_5 (.ZN (n_0_4), .A1 (y), .A2 (n_0_1), .A3 (n_0_3));
AND2_X1 i_0_3 (.ZN (n_0_3), .A1 (cin), .A2 (x));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (cin), .A2 (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_282

module PartialAdder__1_283 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_189 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_192 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_195 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_198 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_201 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_204 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_207 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_210 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_213 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_216 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_219 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_222 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_225 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_228 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_231 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_234 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_237 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_240 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_243 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_246 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_249 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_252 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_255 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_258 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_261 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_264 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_267 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_270 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_273 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_276 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_279 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_282 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_283

module halfAdder__1_92 (x, y, sum, cout);

output cout;
output sum;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //halfAdder__1_92

module fullAdder__1_95 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_95

module fullAdder__1_98 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_98

module fullAdder__1_101 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_101

module fullAdder__1_104 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_104

module fullAdder__1_107 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_107

module fullAdder__1_110 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_110

module fullAdder__1_113 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_113

module fullAdder__1_116 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_116

module fullAdder__1_119 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_119

module fullAdder__1_122 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_122

module fullAdder__1_125 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_125

module fullAdder__1_128 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_128

module fullAdder__1_131 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_131

module fullAdder__1_134 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_134

module fullAdder__1_137 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_137

module fullAdder__1_140 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_140

module fullAdder__1_143 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_143

module fullAdder__1_146 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_3), .A2 (x), .B1 (n_0_4), .B2 (n_0_1));
INV_X1 i_0_5 (.ZN (n_0_4), .A (x));
INV_X1 i_0_3 (.ZN (n_0_3), .A (n_0_1));
XNOR2_X1 i_0_2 (.ZN (n_0_1), .A (y), .B (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_146

module fullAdder__1_149 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
OR3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (y));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (y), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (y));
NOR2_X1 i_0_1 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (x), .A2 (cin));

endmodule //fullAdder__1_149

module fullAdder__1_152 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NOR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (cin));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //fullAdder__1_152

module fullAdder__1_155 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_155

module fullAdder__1_158 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_7));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (x), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (n_0_4));
INV_X1 i_0_4 (.ZN (sum), .A (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_2), .A (y));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (x), .A2 (cin));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (x), .A2 (cin));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_0), .B2 (n_0_2));

endmodule //fullAdder__1_158

module fullAdder__1_161 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_3), .A (y), .B (cin));
INV_X1 i_0_2 (.ZN (n_0_1), .A (x));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_161

module fullAdder__1_164 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X2 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_164

module fullAdder__1_167 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X1 i_0_6 (.ZN (sum), .A1 (n_0_1), .A2 (n_0_3), .B1 (x), .B2 (n_0_4));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_4 (.ZN (n_0_3), .A (y), .B (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (cin));
INV_X1 i_0_1 (.ZN (n_0_1), .A (x));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (y), .B1 (x), .B2 (cin));

endmodule //fullAdder__1_167

module fullAdder__1_170 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


XNOR2_X1 i_0_9 (.ZN (n_0_7), .A (y), .B (cin));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (x), .A2 (n_0_7));
OAI21_X1 i_0_7 (.ZN (sum), .A (n_0_6), .B1 (x), .B2 (n_0_7));
INV_X1 i_0_6 (.ZN (n_0_5), .A (y));
NOR2_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_3), .A1 (x), .A2 (cin));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_3), .B1 (n_0_4), .B2 (n_0_5));

endmodule //fullAdder__1_170

module fullAdder__1_173 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (x));
XNOR2_X1 i_0_7 (.ZN (n_0_5), .A (y), .B (cin));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_5));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (y), .A2 (cin));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_173

module fullAdder__1_176 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (x));
INV_X1 i_0_9 (.ZN (n_0_7), .A (cin));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (y), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (n_0_6));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_2 (.ZN (sum), .A (n_0_1));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_176

module fullAdder__1_179 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X2 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_179

module fullAdder__1_182 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_2;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (x), .B1 (n_0_1), .B2 (n_0_3));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (x), .A2 (n_0_1), .A3 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_3), .A1 (y), .A2 (cin));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (y), .A2 (cin));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__1_182

module fullAdder__1_185 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X1 i_0_7 (.ZN (sum), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (y), .B1 (n_0_3), .B2 (n_0_0));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_3), .A2 (y), .A3 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
OAI21_X1 i_0_3 (.ZN (cout), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_2), .A1 (cin), .A2 (x));
INV_X1 i_0_1 (.ZN (n_0_1), .A (y));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (cin), .A2 (x));

endmodule //fullAdder__1_185

module PartialAdder__1_186 (a, b, c, s1, c1);

output [31:0] c1;
output [32:0] s1;
input [32:0] a;
input [31:0] b;
input [31:0] c;


halfAdder__1_92 ha1 (.cout (c1[0]), .sum (s1[0]), .x (a[1]), .y (b[0]));
fullAdder__1_95 fa1 (.cout (c1[1]), .sum (s1[1]), .cin (c[0]), .x (a[2]), .y (b[1]));
fullAdder__1_98 fa2 (.cout (c1[2]), .sum (s1[2]), .cin (c[1]), .x (a[3]), .y (b[2]));
fullAdder__1_101 fa3 (.cout (c1[3]), .sum (s1[3]), .cin (c[2]), .x (a[4]), .y (b[3]));
fullAdder__1_104 fa4 (.cout (c1[4]), .sum (s1[4]), .cin (c[3]), .x (a[5]), .y (b[4]));
fullAdder__1_107 fa5 (.cout (c1[5]), .sum (s1[5]), .cin (c[4]), .x (a[6]), .y (b[5]));
fullAdder__1_110 fa6 (.cout (c1[6]), .sum (s1[6]), .cin (c[5]), .x (a[7]), .y (b[6]));
fullAdder__1_113 fa7 (.cout (c1[7]), .sum (s1[7]), .cin (c[6]), .x (a[8]), .y (b[7]));
fullAdder__1_116 fa8 (.cout (c1[8]), .sum (s1[8]), .cin (c[7]), .x (a[9]), .y (b[8]));
fullAdder__1_119 fa9 (.cout (c1[9]), .sum (s1[9]), .cin (c[8]), .x (a[10]), .y (b[9]));
fullAdder__1_122 fa10 (.cout (c1[10]), .sum (s1[10]), .cin (c[9]), .x (a[11]), .y (b[10]));
fullAdder__1_125 fa11 (.cout (c1[11]), .sum (s1[11]), .cin (c[10]), .x (a[12]), .y (b[11]));
fullAdder__1_128 fa12 (.cout (c1[12]), .sum (s1[12]), .cin (c[11]), .x (a[13]), .y (b[12]));
fullAdder__1_131 fa13 (.cout (c1[13]), .sum (s1[13]), .cin (c[12]), .x (a[14]), .y (b[13]));
fullAdder__1_134 fa14 (.cout (c1[14]), .sum (s1[14]), .cin (c[13]), .x (a[15]), .y (b[14]));
fullAdder__1_137 fa15 (.cout (c1[15]), .sum (s1[15]), .cin (c[14]), .x (a[16]), .y (b[15]));
fullAdder__1_140 fa16 (.cout (c1[16]), .sum (s1[16]), .cin (c[15]), .x (a[17]), .y (b[16]));
fullAdder__1_143 fa17 (.cout (c1[17]), .sum (s1[17]), .cin (c[16]), .x (a[18]), .y (b[17]));
fullAdder__1_146 fa18 (.cout (c1[18]), .sum (s1[18]), .cin (c[17]), .x (a[19]), .y (b[18]));
fullAdder__1_149 fa19 (.cout (c1[19]), .sum (s1[19]), .cin (c[18]), .x (a[20]), .y (b[19]));
fullAdder__1_152 fa20 (.cout (c1[20]), .sum (s1[20]), .cin (c[19]), .x (a[21]), .y (b[20]));
fullAdder__1_155 fa21 (.cout (c1[21]), .sum (s1[21]), .cin (c[20]), .x (a[22]), .y (b[21]));
fullAdder__1_158 fa22 (.cout (c1[22]), .sum (s1[22]), .cin (c[21]), .x (a[23]), .y (b[22]));
fullAdder__1_161 fa23 (.cout (c1[23]), .sum (s1[23]), .cin (c[22]), .x (a[24]), .y (b[23]));
fullAdder__1_164 fa24 (.cout (c1[24]), .sum (s1[24]), .cin (c[23]), .x (a[25]), .y (b[24]));
fullAdder__1_167 fa25 (.cout (c1[25]), .sum (s1[25]), .cin (c[24]), .x (a[26]), .y (b[25]));
fullAdder__1_170 fa26 (.cout (c1[26]), .sum (s1[26]), .cin (c[25]), .x (a[27]), .y (b[26]));
fullAdder__1_173 fa27 (.cout (c1[27]), .sum (s1[27]), .cin (c[26]), .x (a[28]), .y (b[27]));
fullAdder__1_176 fa28 (.cout (c1[28]), .sum (s1[28]), .cin (c[27]), .x (a[29]), .y (b[28]));
fullAdder__1_179 fa29 (.cout (c1[29]), .sum (s1[29]), .cin (c[28]), .x (a[30]), .y (b[29]));
fullAdder__1_182 fa30 (.cout (c1[30]), .sum (s1[30]), .cin (c[29]), .x (a[31]), .y (b[30]));
fullAdder__1_185 fa31 (.cout (c1[31]), .sum (s1[31]), .cin (c[30]), .x (a[32]), .y (b[31]));

endmodule //PartialAdder__1_186

module TreeMultiplierCirc (a, b, out);

output [63:0] out;
input [31:0] a;
input [31:0] b;
wire \c1[1][31] ;
wire \c1[1][30] ;
wire \c1[1][29] ;
wire \c1[1][28] ;
wire \c1[1][27] ;
wire \c1[1][26] ;
wire \c1[1][25] ;
wire \c1[1][24] ;
wire \c1[1][23] ;
wire \c1[1][22] ;
wire \c1[1][21] ;
wire \c1[1][20] ;
wire \c1[1][19] ;
wire \c1[1][18] ;
wire \c1[1][17] ;
wire \c1[1][16] ;
wire \c1[1][15] ;
wire \c1[1][14] ;
wire \c1[1][13] ;
wire \c1[1][12] ;
wire \c1[1][11] ;
wire \c1[1][10] ;
wire \c1[1][9] ;
wire \c1[1][8] ;
wire \c1[1][7] ;
wire \c1[1][6] ;
wire \c1[1][5] ;
wire \c1[1][4] ;
wire \c1[1][3] ;
wire \c1[1][2] ;
wire \c1[1][1] ;
wire \c1[1][0] ;
wire n_39_0;
wire n_39_1;
wire n_39_2;
wire n_39_3;
wire n_39_4;
wire n_39_5;
wire n_39_6;
wire n_39_7;
wire n_39_8;
wire n_39_9;
wire n_39_10;
wire n_39_11;
wire n_39_12;
wire n_39_13;
wire n_39_14;
wire n_39_15;
wire n_39_16;
wire n_39_17;
wire n_39_18;
wire n_39_19;
wire n_39_20;
wire n_39_21;
wire n_39_22;
wire n_39_23;
wire n_39_24;
wire n_39_25;
wire n_39_26;
wire n_39_27;
wire n_39_28;
wire n_39_29;
wire n_39_30;
wire \c1[2][31] ;
wire \c1[2][30] ;
wire \c1[2][29] ;
wire \c1[2][28] ;
wire \c1[2][27] ;
wire \c1[2][26] ;
wire \c1[2][25] ;
wire \c1[2][24] ;
wire \c1[2][23] ;
wire \c1[2][22] ;
wire \c1[2][21] ;
wire \c1[2][20] ;
wire \c1[2][19] ;
wire \c1[2][18] ;
wire \c1[2][17] ;
wire \c1[2][16] ;
wire \c1[2][15] ;
wire \c1[2][14] ;
wire \c1[2][13] ;
wire \c1[2][12] ;
wire \c1[2][11] ;
wire \c1[2][10] ;
wire \c1[2][9] ;
wire \c1[2][8] ;
wire \c1[2][7] ;
wire \c1[2][6] ;
wire \c1[2][5] ;
wire \c1[2][4] ;
wire \c1[2][3] ;
wire \c1[2][2] ;
wire \c1[2][1] ;
wire \c1[2][0] ;
wire n_39_32;
wire n_39_33;
wire n_39_34;
wire n_39_35;
wire n_39_36;
wire n_39_37;
wire n_39_38;
wire n_39_39;
wire n_39_40;
wire n_39_41;
wire n_39_42;
wire n_39_43;
wire n_39_44;
wire n_39_45;
wire n_39_46;
wire n_39_47;
wire n_39_48;
wire n_39_49;
wire n_39_50;
wire n_39_51;
wire n_39_52;
wire n_39_53;
wire n_39_54;
wire n_39_55;
wire n_39_56;
wire n_39_57;
wire n_39_58;
wire n_39_59;
wire n_39_60;
wire n_39_61;
wire n_39_62;
wire \c1[3][31] ;
wire \c1[3][30] ;
wire \c1[3][29] ;
wire \c1[3][28] ;
wire \c1[3][27] ;
wire \c1[3][26] ;
wire \c1[3][25] ;
wire \c1[3][24] ;
wire \c1[3][23] ;
wire \c1[3][22] ;
wire \c1[3][21] ;
wire \c1[3][20] ;
wire \c1[3][19] ;
wire \c1[3][18] ;
wire \c1[3][17] ;
wire \c1[3][16] ;
wire \c1[3][15] ;
wire \c1[3][14] ;
wire \c1[3][13] ;
wire \c1[3][12] ;
wire \c1[3][11] ;
wire \c1[3][10] ;
wire \c1[3][9] ;
wire \c1[3][8] ;
wire \c1[3][7] ;
wire \c1[3][6] ;
wire \c1[3][5] ;
wire \c1[3][4] ;
wire \c1[3][3] ;
wire \c1[3][2] ;
wire \c1[3][1] ;
wire \c1[3][0] ;
wire n_39_64;
wire n_39_65;
wire n_39_66;
wire n_39_67;
wire n_39_68;
wire n_39_69;
wire n_39_70;
wire n_39_71;
wire n_39_72;
wire n_39_73;
wire n_39_74;
wire n_39_75;
wire n_39_76;
wire n_39_77;
wire n_39_78;
wire n_39_79;
wire n_39_80;
wire n_39_81;
wire n_39_82;
wire n_39_83;
wire n_39_84;
wire n_39_85;
wire n_39_86;
wire n_39_87;
wire n_39_88;
wire n_39_89;
wire n_39_90;
wire n_39_91;
wire n_39_92;
wire n_39_93;
wire n_39_94;
wire \c1[4][31] ;
wire \c1[4][30] ;
wire \c1[4][29] ;
wire \c1[4][28] ;
wire \c1[4][27] ;
wire \c1[4][26] ;
wire \c1[4][25] ;
wire \c1[4][24] ;
wire \c1[4][23] ;
wire \c1[4][22] ;
wire \c1[4][21] ;
wire \c1[4][20] ;
wire \c1[4][19] ;
wire \c1[4][18] ;
wire \c1[4][17] ;
wire \c1[4][16] ;
wire \c1[4][15] ;
wire \c1[4][14] ;
wire \c1[4][13] ;
wire \c1[4][12] ;
wire \c1[4][11] ;
wire \c1[4][10] ;
wire \c1[4][9] ;
wire \c1[4][8] ;
wire \c1[4][7] ;
wire \c1[4][6] ;
wire \c1[4][5] ;
wire \c1[4][4] ;
wire \c1[4][3] ;
wire \c1[4][2] ;
wire \c1[4][1] ;
wire \c1[4][0] ;
wire n_39_96;
wire n_39_97;
wire n_39_98;
wire n_39_99;
wire n_39_100;
wire n_39_101;
wire n_39_102;
wire n_39_103;
wire n_39_104;
wire n_39_105;
wire n_39_106;
wire n_39_107;
wire n_39_108;
wire n_39_109;
wire n_39_110;
wire n_39_111;
wire n_39_112;
wire n_39_113;
wire n_39_114;
wire n_39_115;
wire n_39_116;
wire n_39_117;
wire n_39_118;
wire n_39_119;
wire n_39_120;
wire n_39_121;
wire n_39_122;
wire n_39_123;
wire n_39_124;
wire n_39_125;
wire n_39_126;
wire \c1[5][31] ;
wire \c1[5][30] ;
wire \c1[5][29] ;
wire \c1[5][28] ;
wire \c1[5][27] ;
wire \c1[5][26] ;
wire \c1[5][25] ;
wire \c1[5][24] ;
wire \c1[5][23] ;
wire \c1[5][22] ;
wire \c1[5][21] ;
wire \c1[5][20] ;
wire \c1[5][19] ;
wire \c1[5][18] ;
wire \c1[5][17] ;
wire \c1[5][16] ;
wire \c1[5][15] ;
wire \c1[5][14] ;
wire \c1[5][13] ;
wire \c1[5][12] ;
wire \c1[5][11] ;
wire \c1[5][10] ;
wire \c1[5][9] ;
wire \c1[5][8] ;
wire \c1[5][7] ;
wire \c1[5][6] ;
wire \c1[5][5] ;
wire \c1[5][4] ;
wire \c1[5][3] ;
wire \c1[5][2] ;
wire \c1[5][1] ;
wire \c1[5][0] ;
wire n_39_128;
wire n_39_129;
wire n_39_130;
wire n_39_131;
wire n_39_132;
wire n_39_133;
wire n_39_134;
wire n_39_135;
wire n_39_136;
wire n_39_137;
wire n_39_138;
wire n_39_139;
wire n_39_140;
wire n_39_141;
wire n_39_142;
wire n_39_143;
wire n_39_144;
wire n_39_145;
wire n_39_146;
wire n_39_147;
wire n_39_148;
wire n_39_149;
wire n_39_150;
wire n_39_151;
wire n_39_152;
wire n_39_153;
wire n_39_154;
wire n_39_155;
wire n_39_156;
wire n_39_157;
wire n_39_158;
wire \c1[6][31] ;
wire \c1[6][30] ;
wire \c1[6][29] ;
wire \c1[6][28] ;
wire \c1[6][27] ;
wire \c1[6][26] ;
wire \c1[6][25] ;
wire \c1[6][24] ;
wire \c1[6][23] ;
wire \c1[6][22] ;
wire \c1[6][21] ;
wire \c1[6][20] ;
wire \c1[6][19] ;
wire \c1[6][18] ;
wire \c1[6][17] ;
wire \c1[6][16] ;
wire \c1[6][15] ;
wire \c1[6][14] ;
wire \c1[6][13] ;
wire \c1[6][12] ;
wire \c1[6][11] ;
wire \c1[6][10] ;
wire \c1[6][9] ;
wire \c1[6][8] ;
wire \c1[6][7] ;
wire \c1[6][6] ;
wire \c1[6][5] ;
wire \c1[6][4] ;
wire \c1[6][3] ;
wire \c1[6][2] ;
wire \c1[6][1] ;
wire \c1[6][0] ;
wire n_39_160;
wire n_39_161;
wire n_39_162;
wire n_39_163;
wire n_39_164;
wire n_39_165;
wire n_39_166;
wire n_39_167;
wire n_39_168;
wire n_39_169;
wire n_39_170;
wire n_39_171;
wire n_39_172;
wire n_39_173;
wire n_39_174;
wire n_39_175;
wire n_39_176;
wire n_39_177;
wire n_39_178;
wire n_39_179;
wire n_39_180;
wire n_39_181;
wire n_39_182;
wire n_39_183;
wire n_39_184;
wire n_39_185;
wire n_39_186;
wire n_39_187;
wire n_39_188;
wire n_39_189;
wire n_39_190;
wire \c1[7][31] ;
wire \c1[7][30] ;
wire \c1[7][29] ;
wire \c1[7][28] ;
wire \c1[7][27] ;
wire \c1[7][26] ;
wire \c1[7][25] ;
wire \c1[7][24] ;
wire \c1[7][23] ;
wire \c1[7][22] ;
wire \c1[7][21] ;
wire \c1[7][20] ;
wire \c1[7][19] ;
wire \c1[7][18] ;
wire \c1[7][17] ;
wire \c1[7][16] ;
wire \c1[7][15] ;
wire \c1[7][14] ;
wire \c1[7][13] ;
wire \c1[7][12] ;
wire \c1[7][11] ;
wire \c1[7][10] ;
wire \c1[7][9] ;
wire \c1[7][8] ;
wire \c1[7][7] ;
wire \c1[7][6] ;
wire \c1[7][5] ;
wire \c1[7][4] ;
wire \c1[7][3] ;
wire \c1[7][2] ;
wire \c1[7][1] ;
wire \c1[7][0] ;
wire n_39_192;
wire n_39_193;
wire n_39_194;
wire n_39_195;
wire n_39_196;
wire n_39_197;
wire n_39_198;
wire n_39_199;
wire n_39_200;
wire n_39_201;
wire n_39_202;
wire n_39_203;
wire n_39_204;
wire n_39_205;
wire n_39_206;
wire n_39_207;
wire n_39_208;
wire n_39_209;
wire n_39_210;
wire n_39_211;
wire n_39_212;
wire n_39_213;
wire n_39_214;
wire n_39_215;
wire n_39_216;
wire n_39_217;
wire n_39_218;
wire n_39_219;
wire n_39_220;
wire n_39_221;
wire n_39_222;
wire \c1[8][31] ;
wire \c1[8][30] ;
wire \c1[8][29] ;
wire \c1[8][28] ;
wire \c1[8][27] ;
wire \c1[8][26] ;
wire \c1[8][25] ;
wire \c1[8][24] ;
wire \c1[8][23] ;
wire \c1[8][22] ;
wire \c1[8][21] ;
wire \c1[8][20] ;
wire \c1[8][19] ;
wire \c1[8][18] ;
wire \c1[8][17] ;
wire \c1[8][16] ;
wire \c1[8][15] ;
wire \c1[8][14] ;
wire \c1[8][13] ;
wire \c1[8][12] ;
wire \c1[8][11] ;
wire \c1[8][10] ;
wire \c1[8][9] ;
wire \c1[8][8] ;
wire \c1[8][7] ;
wire \c1[8][6] ;
wire \c1[8][5] ;
wire \c1[8][4] ;
wire \c1[8][3] ;
wire \c1[8][2] ;
wire \c1[8][1] ;
wire \c1[8][0] ;
wire n_39_224;
wire n_39_225;
wire n_39_226;
wire n_39_227;
wire n_39_228;
wire n_39_229;
wire n_39_230;
wire n_39_231;
wire n_39_232;
wire n_39_233;
wire n_39_234;
wire n_39_235;
wire n_39_236;
wire n_39_237;
wire n_39_238;
wire n_39_239;
wire n_39_240;
wire n_39_241;
wire n_39_242;
wire n_39_243;
wire n_39_244;
wire n_39_245;
wire n_39_246;
wire n_39_247;
wire n_39_248;
wire n_39_249;
wire n_39_250;
wire n_39_251;
wire n_39_252;
wire n_39_253;
wire n_39_254;
wire \c1[9][31] ;
wire \c1[9][30] ;
wire \c1[9][29] ;
wire \c1[9][28] ;
wire \c1[9][27] ;
wire \c1[9][26] ;
wire \c1[9][25] ;
wire \c1[9][24] ;
wire \c1[9][23] ;
wire \c1[9][22] ;
wire \c1[9][21] ;
wire \c1[9][20] ;
wire \c1[9][19] ;
wire \c1[9][18] ;
wire \c1[9][17] ;
wire \c1[9][16] ;
wire \c1[9][15] ;
wire \c1[9][14] ;
wire \c1[9][13] ;
wire \c1[9][12] ;
wire \c1[9][11] ;
wire \c1[9][10] ;
wire \c1[9][9] ;
wire \c1[9][8] ;
wire \c1[9][7] ;
wire \c1[9][6] ;
wire \c1[9][5] ;
wire \c1[9][4] ;
wire \c1[9][3] ;
wire \c1[9][2] ;
wire \c1[9][1] ;
wire \c1[9][0] ;
wire n_39_256;
wire n_39_257;
wire n_39_258;
wire n_39_259;
wire n_39_260;
wire n_39_261;
wire n_39_262;
wire n_39_263;
wire n_39_264;
wire n_39_265;
wire n_39_266;
wire n_39_267;
wire n_39_268;
wire n_39_269;
wire n_39_270;
wire n_39_271;
wire n_39_272;
wire n_39_273;
wire n_39_274;
wire n_39_275;
wire n_39_276;
wire n_39_277;
wire n_39_278;
wire n_39_279;
wire n_39_280;
wire n_39_281;
wire n_39_282;
wire n_39_283;
wire n_39_284;
wire n_39_285;
wire n_39_286;
wire \c1[10][31] ;
wire \c1[10][30] ;
wire \c1[10][29] ;
wire \c1[10][28] ;
wire \c1[10][27] ;
wire \c1[10][26] ;
wire \c1[10][25] ;
wire \c1[10][24] ;
wire \c1[10][23] ;
wire \c1[10][22] ;
wire \c1[10][21] ;
wire \c1[10][20] ;
wire \c1[10][19] ;
wire \c1[10][18] ;
wire \c1[10][17] ;
wire \c1[10][16] ;
wire \c1[10][15] ;
wire \c1[10][14] ;
wire \c1[10][13] ;
wire \c1[10][12] ;
wire \c1[10][11] ;
wire \c1[10][10] ;
wire \c1[10][9] ;
wire \c1[10][8] ;
wire \c1[10][7] ;
wire \c1[10][6] ;
wire \c1[10][5] ;
wire \c1[10][4] ;
wire \c1[10][3] ;
wire \c1[10][2] ;
wire \c1[10][1] ;
wire \c1[10][0] ;
wire n_39_288;
wire n_39_289;
wire n_39_290;
wire n_39_291;
wire n_39_292;
wire n_39_293;
wire n_39_294;
wire n_39_295;
wire n_39_296;
wire n_39_297;
wire n_39_298;
wire n_39_299;
wire n_39_300;
wire n_39_301;
wire n_39_302;
wire n_39_303;
wire n_39_304;
wire n_39_305;
wire n_39_306;
wire n_39_307;
wire n_39_308;
wire n_39_309;
wire n_39_310;
wire n_39_311;
wire n_39_312;
wire n_39_313;
wire n_39_314;
wire n_39_315;
wire n_39_316;
wire n_39_317;
wire n_39_318;
wire \c1[11][31] ;
wire \c1[11][30] ;
wire \c1[11][29] ;
wire \c1[11][28] ;
wire \c1[11][27] ;
wire \c1[11][26] ;
wire \c1[11][25] ;
wire \c1[11][24] ;
wire \c1[11][23] ;
wire \c1[11][22] ;
wire \c1[11][21] ;
wire \c1[11][20] ;
wire \c1[11][19] ;
wire \c1[11][18] ;
wire \c1[11][17] ;
wire \c1[11][16] ;
wire \c1[11][15] ;
wire \c1[11][14] ;
wire \c1[11][13] ;
wire \c1[11][12] ;
wire \c1[11][11] ;
wire \c1[11][10] ;
wire \c1[11][9] ;
wire \c1[11][8] ;
wire \c1[11][7] ;
wire \c1[11][6] ;
wire \c1[11][5] ;
wire \c1[11][4] ;
wire \c1[11][3] ;
wire \c1[11][2] ;
wire \c1[11][1] ;
wire \c1[11][0] ;
wire n_39_320;
wire n_39_321;
wire n_39_322;
wire n_39_323;
wire n_39_324;
wire n_39_325;
wire n_39_326;
wire n_39_327;
wire n_39_328;
wire n_39_329;
wire n_39_330;
wire n_39_331;
wire n_39_332;
wire n_39_333;
wire n_39_334;
wire n_39_335;
wire n_39_336;
wire n_39_337;
wire n_39_338;
wire n_39_339;
wire n_39_340;
wire n_39_341;
wire n_39_342;
wire n_39_343;
wire n_39_344;
wire n_39_345;
wire n_39_346;
wire n_39_347;
wire n_39_348;
wire n_39_349;
wire n_39_350;
wire \c1[12][31] ;
wire \c1[12][30] ;
wire \c1[12][29] ;
wire \c1[12][28] ;
wire \c1[12][27] ;
wire \c1[12][26] ;
wire \c1[12][25] ;
wire \c1[12][24] ;
wire \c1[12][23] ;
wire \c1[12][22] ;
wire \c1[12][21] ;
wire \c1[12][20] ;
wire \c1[12][19] ;
wire \c1[12][18] ;
wire \c1[12][17] ;
wire \c1[12][16] ;
wire \c1[12][15] ;
wire \c1[12][14] ;
wire \c1[12][13] ;
wire \c1[12][12] ;
wire \c1[12][11] ;
wire \c1[12][10] ;
wire \c1[12][9] ;
wire \c1[12][8] ;
wire \c1[12][7] ;
wire \c1[12][6] ;
wire \c1[12][5] ;
wire \c1[12][4] ;
wire \c1[12][3] ;
wire \c1[12][2] ;
wire \c1[12][1] ;
wire \c1[12][0] ;
wire n_39_352;
wire n_39_353;
wire n_39_354;
wire n_39_355;
wire n_39_356;
wire n_39_357;
wire n_39_358;
wire n_39_359;
wire n_39_360;
wire n_39_361;
wire n_39_362;
wire n_39_363;
wire n_39_364;
wire n_39_365;
wire n_39_366;
wire n_39_367;
wire n_39_368;
wire n_39_369;
wire n_39_370;
wire n_39_371;
wire n_39_372;
wire n_39_373;
wire n_39_374;
wire n_39_375;
wire n_39_376;
wire n_39_377;
wire n_39_378;
wire n_39_379;
wire n_39_380;
wire n_39_381;
wire n_39_382;
wire \c1[13][31] ;
wire \c1[13][30] ;
wire \c1[13][29] ;
wire \c1[13][28] ;
wire \c1[13][27] ;
wire \c1[13][26] ;
wire \c1[13][25] ;
wire \c1[13][24] ;
wire \c1[13][23] ;
wire \c1[13][22] ;
wire \c1[13][21] ;
wire \c1[13][20] ;
wire \c1[13][19] ;
wire \c1[13][18] ;
wire \c1[13][17] ;
wire \c1[13][16] ;
wire \c1[13][15] ;
wire \c1[13][14] ;
wire \c1[13][13] ;
wire \c1[13][12] ;
wire \c1[13][11] ;
wire \c1[13][10] ;
wire \c1[13][9] ;
wire \c1[13][8] ;
wire \c1[13][7] ;
wire \c1[13][6] ;
wire \c1[13][5] ;
wire \c1[13][4] ;
wire \c1[13][3] ;
wire \c1[13][2] ;
wire \c1[13][1] ;
wire \c1[13][0] ;
wire n_39_384;
wire n_39_385;
wire n_39_386;
wire n_39_387;
wire n_39_388;
wire n_39_389;
wire n_39_390;
wire n_39_391;
wire n_39_392;
wire n_39_393;
wire n_39_394;
wire n_39_395;
wire n_39_396;
wire n_39_397;
wire n_39_398;
wire n_39_399;
wire n_39_400;
wire n_39_401;
wire n_39_402;
wire n_39_403;
wire n_39_404;
wire n_39_405;
wire n_39_406;
wire n_39_407;
wire n_39_408;
wire n_39_409;
wire n_39_410;
wire n_39_411;
wire n_39_412;
wire n_39_413;
wire n_39_414;
wire \c1[14][31] ;
wire \c1[14][30] ;
wire \c1[14][29] ;
wire \c1[14][28] ;
wire \c1[14][27] ;
wire \c1[14][26] ;
wire \c1[14][25] ;
wire \c1[14][24] ;
wire \c1[14][23] ;
wire \c1[14][22] ;
wire \c1[14][21] ;
wire \c1[14][20] ;
wire \c1[14][19] ;
wire \c1[14][18] ;
wire \c1[14][17] ;
wire \c1[14][16] ;
wire \c1[14][15] ;
wire \c1[14][14] ;
wire \c1[14][13] ;
wire \c1[14][12] ;
wire \c1[14][11] ;
wire \c1[14][10] ;
wire \c1[14][9] ;
wire \c1[14][8] ;
wire \c1[14][7] ;
wire \c1[14][6] ;
wire \c1[14][5] ;
wire \c1[14][4] ;
wire \c1[14][3] ;
wire \c1[14][2] ;
wire \c1[14][1] ;
wire \c1[14][0] ;
wire n_39_416;
wire n_39_417;
wire n_39_418;
wire n_39_419;
wire n_39_420;
wire n_39_421;
wire n_39_422;
wire n_39_423;
wire n_39_424;
wire n_39_425;
wire n_39_426;
wire n_39_427;
wire n_39_428;
wire n_39_429;
wire n_39_430;
wire n_39_431;
wire n_39_432;
wire n_39_433;
wire n_39_434;
wire n_39_435;
wire n_39_436;
wire n_39_437;
wire n_39_438;
wire n_39_439;
wire n_39_440;
wire n_39_441;
wire n_39_442;
wire n_39_443;
wire n_39_444;
wire n_39_445;
wire n_39_446;
wire \c1[15][31] ;
wire \c1[15][30] ;
wire \c1[15][29] ;
wire \c1[15][28] ;
wire \c1[15][27] ;
wire \c1[15][26] ;
wire \c1[15][25] ;
wire \c1[15][24] ;
wire \c1[15][23] ;
wire \c1[15][22] ;
wire \c1[15][21] ;
wire \c1[15][20] ;
wire \c1[15][19] ;
wire \c1[15][18] ;
wire \c1[15][17] ;
wire \c1[15][16] ;
wire \c1[15][15] ;
wire \c1[15][14] ;
wire \c1[15][13] ;
wire \c1[15][12] ;
wire \c1[15][11] ;
wire \c1[15][10] ;
wire \c1[15][9] ;
wire \c1[15][8] ;
wire \c1[15][7] ;
wire \c1[15][6] ;
wire \c1[15][5] ;
wire \c1[15][4] ;
wire \c1[15][3] ;
wire \c1[15][2] ;
wire \c1[15][1] ;
wire \c1[15][0] ;
wire n_39_448;
wire n_39_449;
wire n_39_450;
wire n_39_451;
wire n_39_452;
wire n_39_453;
wire n_39_454;
wire n_39_455;
wire n_39_456;
wire n_39_457;
wire n_39_458;
wire n_39_459;
wire n_39_460;
wire n_39_461;
wire n_39_462;
wire n_39_463;
wire n_39_464;
wire n_39_465;
wire n_39_466;
wire n_39_467;
wire n_39_468;
wire n_39_469;
wire n_39_470;
wire n_39_471;
wire n_39_472;
wire n_39_473;
wire n_39_474;
wire n_39_475;
wire n_39_476;
wire n_39_477;
wire n_39_478;
wire \c1[16][31] ;
wire \c1[16][30] ;
wire \c1[16][29] ;
wire \c1[16][28] ;
wire \c1[16][27] ;
wire \c1[16][26] ;
wire \c1[16][25] ;
wire \c1[16][24] ;
wire \c1[16][23] ;
wire \c1[16][22] ;
wire \c1[16][21] ;
wire \c1[16][20] ;
wire \c1[16][19] ;
wire \c1[16][18] ;
wire \c1[16][17] ;
wire \c1[16][16] ;
wire \c1[16][15] ;
wire \c1[16][14] ;
wire \c1[16][13] ;
wire \c1[16][12] ;
wire \c1[16][11] ;
wire \c1[16][10] ;
wire \c1[16][9] ;
wire \c1[16][8] ;
wire \c1[16][7] ;
wire \c1[16][6] ;
wire \c1[16][5] ;
wire \c1[16][4] ;
wire \c1[16][3] ;
wire \c1[16][2] ;
wire \c1[16][1] ;
wire \c1[16][0] ;
wire n_39_480;
wire n_39_481;
wire n_39_482;
wire n_39_483;
wire n_39_484;
wire n_39_485;
wire n_39_486;
wire n_39_487;
wire n_39_488;
wire n_39_489;
wire n_39_490;
wire n_39_491;
wire n_39_492;
wire n_39_493;
wire n_39_494;
wire n_39_495;
wire n_39_496;
wire n_39_497;
wire n_39_498;
wire n_39_499;
wire n_39_500;
wire n_39_501;
wire n_39_502;
wire n_39_503;
wire n_39_504;
wire n_39_505;
wire n_39_506;
wire n_39_507;
wire n_39_508;
wire n_39_509;
wire n_39_510;
wire \c1[17][31] ;
wire \c1[17][30] ;
wire \c1[17][29] ;
wire \c1[17][28] ;
wire \c1[17][27] ;
wire \c1[17][26] ;
wire \c1[17][25] ;
wire \c1[17][24] ;
wire \c1[17][23] ;
wire \c1[17][22] ;
wire \c1[17][21] ;
wire \c1[17][20] ;
wire \c1[17][19] ;
wire \c1[17][18] ;
wire \c1[17][17] ;
wire \c1[17][16] ;
wire \c1[17][15] ;
wire \c1[17][14] ;
wire \c1[17][13] ;
wire \c1[17][12] ;
wire \c1[17][11] ;
wire \c1[17][10] ;
wire \c1[17][9] ;
wire \c1[17][8] ;
wire \c1[17][7] ;
wire \c1[17][6] ;
wire \c1[17][5] ;
wire \c1[17][4] ;
wire \c1[17][3] ;
wire \c1[17][2] ;
wire \c1[17][1] ;
wire \c1[17][0] ;
wire n_39_512;
wire n_39_513;
wire n_39_514;
wire n_39_515;
wire n_39_516;
wire n_39_517;
wire n_39_518;
wire n_39_519;
wire n_39_520;
wire n_39_521;
wire n_39_522;
wire n_39_523;
wire n_39_524;
wire n_39_525;
wire n_39_526;
wire n_39_527;
wire n_39_528;
wire n_39_529;
wire n_39_530;
wire n_39_531;
wire n_39_532;
wire n_39_533;
wire n_39_534;
wire n_39_535;
wire n_39_536;
wire n_39_537;
wire n_39_538;
wire n_39_539;
wire n_39_540;
wire n_39_541;
wire n_39_542;
wire \c1[18][31] ;
wire \c1[18][30] ;
wire \c1[18][29] ;
wire \c1[18][28] ;
wire \c1[18][27] ;
wire \c1[18][26] ;
wire \c1[18][25] ;
wire \c1[18][24] ;
wire \c1[18][23] ;
wire \c1[18][22] ;
wire \c1[18][21] ;
wire \c1[18][20] ;
wire \c1[18][19] ;
wire \c1[18][18] ;
wire \c1[18][17] ;
wire \c1[18][16] ;
wire \c1[18][15] ;
wire \c1[18][14] ;
wire \c1[18][13] ;
wire \c1[18][12] ;
wire \c1[18][11] ;
wire \c1[18][10] ;
wire \c1[18][9] ;
wire \c1[18][8] ;
wire \c1[18][7] ;
wire \c1[18][6] ;
wire \c1[18][5] ;
wire \c1[18][4] ;
wire \c1[18][3] ;
wire \c1[18][2] ;
wire \c1[18][1] ;
wire \c1[18][0] ;
wire n_39_544;
wire n_39_545;
wire n_39_546;
wire n_39_547;
wire n_39_548;
wire n_39_549;
wire n_39_550;
wire n_39_551;
wire n_39_552;
wire n_39_553;
wire n_39_554;
wire n_39_555;
wire n_39_556;
wire n_39_557;
wire n_39_558;
wire n_39_559;
wire n_39_560;
wire n_39_561;
wire n_39_562;
wire n_39_563;
wire n_39_564;
wire n_39_565;
wire n_39_566;
wire n_39_567;
wire n_39_568;
wire n_39_569;
wire n_39_570;
wire n_39_571;
wire n_39_572;
wire n_39_573;
wire n_39_574;
wire \c1[19][31] ;
wire \c1[19][30] ;
wire \c1[19][29] ;
wire \c1[19][28] ;
wire \c1[19][27] ;
wire \c1[19][26] ;
wire \c1[19][25] ;
wire \c1[19][24] ;
wire \c1[19][23] ;
wire \c1[19][22] ;
wire \c1[19][21] ;
wire \c1[19][20] ;
wire \c1[19][19] ;
wire \c1[19][18] ;
wire \c1[19][17] ;
wire \c1[19][16] ;
wire \c1[19][15] ;
wire \c1[19][14] ;
wire \c1[19][13] ;
wire \c1[19][12] ;
wire \c1[19][11] ;
wire \c1[19][10] ;
wire \c1[19][9] ;
wire \c1[19][8] ;
wire \c1[19][7] ;
wire \c1[19][6] ;
wire \c1[19][5] ;
wire \c1[19][4] ;
wire \c1[19][3] ;
wire \c1[19][2] ;
wire \c1[19][1] ;
wire \c1[19][0] ;
wire n_39_576;
wire n_39_577;
wire n_39_578;
wire n_39_579;
wire n_39_580;
wire n_39_581;
wire n_39_582;
wire n_39_583;
wire n_39_584;
wire n_39_585;
wire n_39_586;
wire n_39_587;
wire n_39_588;
wire n_39_589;
wire n_39_590;
wire n_39_591;
wire n_39_592;
wire n_39_593;
wire n_39_594;
wire n_39_595;
wire n_39_596;
wire n_39_597;
wire n_39_598;
wire n_39_599;
wire n_39_600;
wire n_39_601;
wire n_39_602;
wire n_39_603;
wire n_39_604;
wire n_39_605;
wire n_39_606;
wire \c1[20][31] ;
wire \c1[20][30] ;
wire \c1[20][29] ;
wire \c1[20][28] ;
wire \c1[20][27] ;
wire \c1[20][26] ;
wire \c1[20][25] ;
wire \c1[20][24] ;
wire \c1[20][23] ;
wire \c1[20][22] ;
wire \c1[20][21] ;
wire \c1[20][20] ;
wire \c1[20][19] ;
wire \c1[20][18] ;
wire \c1[20][17] ;
wire \c1[20][16] ;
wire \c1[20][15] ;
wire \c1[20][14] ;
wire \c1[20][13] ;
wire \c1[20][12] ;
wire \c1[20][11] ;
wire \c1[20][10] ;
wire \c1[20][9] ;
wire \c1[20][8] ;
wire \c1[20][7] ;
wire \c1[20][6] ;
wire \c1[20][5] ;
wire \c1[20][4] ;
wire \c1[20][3] ;
wire \c1[20][2] ;
wire \c1[20][1] ;
wire \c1[20][0] ;
wire n_39_608;
wire n_39_609;
wire n_39_610;
wire n_39_611;
wire n_39_612;
wire n_39_613;
wire n_39_614;
wire n_39_615;
wire n_39_616;
wire n_39_617;
wire n_39_618;
wire n_39_619;
wire n_39_620;
wire n_39_621;
wire n_39_622;
wire n_39_623;
wire n_39_624;
wire n_39_625;
wire n_39_626;
wire n_39_627;
wire n_39_628;
wire n_39_629;
wire n_39_630;
wire n_39_631;
wire n_39_632;
wire n_39_633;
wire n_39_634;
wire n_39_635;
wire n_39_636;
wire n_39_637;
wire n_39_638;
wire \c1[21][31] ;
wire \c1[21][30] ;
wire \c1[21][29] ;
wire \c1[21][28] ;
wire \c1[21][27] ;
wire \c1[21][26] ;
wire \c1[21][25] ;
wire \c1[21][24] ;
wire \c1[21][23] ;
wire \c1[21][22] ;
wire \c1[21][21] ;
wire \c1[21][20] ;
wire \c1[21][19] ;
wire \c1[21][18] ;
wire \c1[21][17] ;
wire \c1[21][16] ;
wire \c1[21][15] ;
wire \c1[21][14] ;
wire \c1[21][13] ;
wire \c1[21][12] ;
wire \c1[21][11] ;
wire \c1[21][10] ;
wire \c1[21][9] ;
wire \c1[21][8] ;
wire \c1[21][7] ;
wire \c1[21][6] ;
wire \c1[21][5] ;
wire \c1[21][4] ;
wire \c1[21][3] ;
wire \c1[21][2] ;
wire \c1[21][1] ;
wire \c1[21][0] ;
wire n_39_640;
wire n_39_641;
wire n_39_642;
wire n_39_643;
wire n_39_644;
wire n_39_645;
wire n_39_646;
wire n_39_647;
wire n_39_648;
wire n_39_649;
wire n_39_650;
wire n_39_651;
wire n_39_652;
wire n_39_653;
wire n_39_654;
wire n_39_655;
wire n_39_656;
wire n_39_657;
wire n_39_658;
wire n_39_659;
wire n_39_660;
wire n_39_661;
wire n_39_662;
wire n_39_663;
wire n_39_664;
wire n_39_665;
wire n_39_666;
wire n_39_667;
wire n_39_668;
wire n_39_669;
wire n_39_670;
wire \c1[22][31] ;
wire \c1[22][30] ;
wire \c1[22][29] ;
wire \c1[22][28] ;
wire \c1[22][27] ;
wire \c1[22][26] ;
wire \c1[22][25] ;
wire \c1[22][24] ;
wire \c1[22][23] ;
wire \c1[22][22] ;
wire \c1[22][21] ;
wire \c1[22][20] ;
wire \c1[22][19] ;
wire \c1[22][18] ;
wire \c1[22][17] ;
wire \c1[22][16] ;
wire \c1[22][15] ;
wire \c1[22][14] ;
wire \c1[22][13] ;
wire \c1[22][12] ;
wire \c1[22][11] ;
wire \c1[22][10] ;
wire \c1[22][9] ;
wire \c1[22][8] ;
wire \c1[22][7] ;
wire \c1[22][6] ;
wire \c1[22][5] ;
wire \c1[22][4] ;
wire \c1[22][3] ;
wire \c1[22][2] ;
wire \c1[22][1] ;
wire \c1[22][0] ;
wire n_39_672;
wire n_39_673;
wire n_39_674;
wire n_39_675;
wire n_39_676;
wire n_39_677;
wire n_39_678;
wire n_39_679;
wire n_39_680;
wire n_39_681;
wire n_39_682;
wire n_39_683;
wire n_39_684;
wire n_39_685;
wire n_39_686;
wire n_39_687;
wire n_39_688;
wire n_39_689;
wire n_39_690;
wire n_39_691;
wire n_39_692;
wire n_39_693;
wire n_39_694;
wire n_39_695;
wire n_39_696;
wire n_39_697;
wire n_39_698;
wire n_39_699;
wire n_39_700;
wire n_39_701;
wire n_39_702;
wire \c1[23][31] ;
wire \c1[23][30] ;
wire \c1[23][29] ;
wire \c1[23][28] ;
wire \c1[23][27] ;
wire \c1[23][26] ;
wire \c1[23][25] ;
wire \c1[23][24] ;
wire \c1[23][23] ;
wire \c1[23][22] ;
wire \c1[23][21] ;
wire \c1[23][20] ;
wire \c1[23][19] ;
wire \c1[23][18] ;
wire \c1[23][17] ;
wire \c1[23][16] ;
wire \c1[23][15] ;
wire \c1[23][14] ;
wire \c1[23][13] ;
wire \c1[23][12] ;
wire \c1[23][11] ;
wire \c1[23][10] ;
wire \c1[23][9] ;
wire \c1[23][8] ;
wire \c1[23][7] ;
wire \c1[23][6] ;
wire \c1[23][5] ;
wire \c1[23][4] ;
wire \c1[23][3] ;
wire \c1[23][2] ;
wire \c1[23][1] ;
wire \c1[23][0] ;
wire n_39_704;
wire n_39_705;
wire n_39_706;
wire n_39_707;
wire n_39_708;
wire n_39_709;
wire n_39_710;
wire n_39_711;
wire n_39_712;
wire n_39_713;
wire n_39_714;
wire n_39_715;
wire n_39_716;
wire n_39_717;
wire n_39_718;
wire n_39_719;
wire n_39_720;
wire n_39_721;
wire n_39_722;
wire n_39_723;
wire n_39_724;
wire n_39_725;
wire n_39_726;
wire n_39_727;
wire n_39_728;
wire n_39_729;
wire n_39_730;
wire n_39_731;
wire n_39_732;
wire n_39_733;
wire n_39_734;
wire \c1[24][31] ;
wire \c1[24][30] ;
wire \c1[24][29] ;
wire \c1[24][28] ;
wire \c1[24][27] ;
wire \c1[24][26] ;
wire \c1[24][25] ;
wire \c1[24][24] ;
wire \c1[24][23] ;
wire \c1[24][22] ;
wire \c1[24][21] ;
wire \c1[24][20] ;
wire \c1[24][19] ;
wire \c1[24][18] ;
wire \c1[24][17] ;
wire \c1[24][16] ;
wire \c1[24][15] ;
wire \c1[24][14] ;
wire \c1[24][13] ;
wire \c1[24][12] ;
wire \c1[24][11] ;
wire \c1[24][10] ;
wire \c1[24][9] ;
wire \c1[24][8] ;
wire \c1[24][7] ;
wire \c1[24][6] ;
wire \c1[24][5] ;
wire \c1[24][4] ;
wire \c1[24][3] ;
wire \c1[24][2] ;
wire \c1[24][1] ;
wire \c1[24][0] ;
wire n_39_736;
wire n_39_737;
wire n_39_738;
wire n_39_739;
wire n_39_740;
wire n_39_741;
wire n_39_742;
wire n_39_743;
wire n_39_744;
wire n_39_745;
wire n_39_746;
wire n_39_747;
wire n_39_748;
wire n_39_749;
wire n_39_750;
wire n_39_751;
wire n_39_752;
wire n_39_753;
wire n_39_754;
wire n_39_755;
wire n_39_756;
wire n_39_757;
wire n_39_758;
wire n_39_759;
wire n_39_760;
wire n_39_761;
wire n_39_762;
wire n_39_763;
wire n_39_764;
wire n_39_765;
wire n_39_766;
wire \c1[25][31] ;
wire \c1[25][30] ;
wire \c1[25][29] ;
wire \c1[25][28] ;
wire \c1[25][27] ;
wire \c1[25][26] ;
wire \c1[25][25] ;
wire \c1[25][24] ;
wire \c1[25][23] ;
wire \c1[25][22] ;
wire \c1[25][21] ;
wire \c1[25][20] ;
wire \c1[25][19] ;
wire \c1[25][18] ;
wire \c1[25][17] ;
wire \c1[25][16] ;
wire \c1[25][15] ;
wire \c1[25][14] ;
wire \c1[25][13] ;
wire \c1[25][12] ;
wire \c1[25][11] ;
wire \c1[25][10] ;
wire \c1[25][9] ;
wire \c1[25][8] ;
wire \c1[25][7] ;
wire \c1[25][6] ;
wire \c1[25][5] ;
wire \c1[25][4] ;
wire \c1[25][3] ;
wire \c1[25][2] ;
wire \c1[25][1] ;
wire \c1[25][0] ;
wire n_39_768;
wire n_39_769;
wire n_39_770;
wire n_39_771;
wire n_39_772;
wire n_39_773;
wire n_39_774;
wire n_39_775;
wire n_39_776;
wire n_39_777;
wire n_39_778;
wire n_39_779;
wire n_39_780;
wire n_39_781;
wire n_39_782;
wire n_39_783;
wire n_39_784;
wire n_39_785;
wire n_39_786;
wire n_39_787;
wire n_39_788;
wire n_39_789;
wire n_39_790;
wire n_39_791;
wire n_39_792;
wire n_39_793;
wire n_39_794;
wire n_39_795;
wire n_39_796;
wire n_39_797;
wire n_39_798;
wire \c1[26][31] ;
wire \c1[26][30] ;
wire \c1[26][29] ;
wire \c1[26][28] ;
wire \c1[26][27] ;
wire \c1[26][26] ;
wire \c1[26][25] ;
wire \c1[26][24] ;
wire \c1[26][23] ;
wire \c1[26][22] ;
wire \c1[26][21] ;
wire \c1[26][20] ;
wire \c1[26][19] ;
wire \c1[26][18] ;
wire \c1[26][17] ;
wire \c1[26][16] ;
wire \c1[26][15] ;
wire \c1[26][14] ;
wire \c1[26][13] ;
wire \c1[26][12] ;
wire \c1[26][11] ;
wire \c1[26][10] ;
wire \c1[26][9] ;
wire \c1[26][8] ;
wire \c1[26][7] ;
wire \c1[26][6] ;
wire \c1[26][5] ;
wire \c1[26][4] ;
wire \c1[26][3] ;
wire \c1[26][2] ;
wire \c1[26][1] ;
wire \c1[26][0] ;
wire n_39_800;
wire n_39_801;
wire n_39_802;
wire n_39_803;
wire n_39_804;
wire n_39_805;
wire n_39_806;
wire n_39_807;
wire n_39_808;
wire n_39_809;
wire n_39_810;
wire n_39_811;
wire n_39_812;
wire n_39_813;
wire n_39_814;
wire n_39_815;
wire n_39_816;
wire n_39_817;
wire n_39_818;
wire n_39_819;
wire n_39_820;
wire n_39_821;
wire n_39_822;
wire n_39_823;
wire n_39_824;
wire n_39_825;
wire n_39_826;
wire n_39_827;
wire n_39_828;
wire n_39_829;
wire n_39_830;
wire \c1[27][31] ;
wire \c1[27][30] ;
wire \c1[27][29] ;
wire \c1[27][28] ;
wire \c1[27][27] ;
wire \c1[27][26] ;
wire \c1[27][25] ;
wire \c1[27][24] ;
wire \c1[27][23] ;
wire \c1[27][22] ;
wire \c1[27][21] ;
wire \c1[27][20] ;
wire \c1[27][19] ;
wire \c1[27][18] ;
wire \c1[27][17] ;
wire \c1[27][16] ;
wire \c1[27][15] ;
wire \c1[27][14] ;
wire \c1[27][13] ;
wire \c1[27][12] ;
wire \c1[27][11] ;
wire \c1[27][10] ;
wire \c1[27][9] ;
wire \c1[27][8] ;
wire \c1[27][7] ;
wire \c1[27][6] ;
wire \c1[27][5] ;
wire \c1[27][4] ;
wire \c1[27][3] ;
wire \c1[27][2] ;
wire \c1[27][1] ;
wire \c1[27][0] ;
wire n_39_832;
wire n_39_833;
wire n_39_834;
wire n_39_835;
wire n_39_836;
wire n_39_837;
wire n_39_838;
wire n_39_839;
wire n_39_840;
wire n_39_841;
wire n_39_842;
wire n_39_843;
wire n_39_844;
wire n_39_845;
wire n_39_846;
wire n_39_847;
wire n_39_848;
wire n_39_849;
wire n_39_850;
wire n_39_851;
wire n_39_852;
wire n_39_853;
wire n_39_854;
wire n_39_855;
wire n_39_856;
wire n_39_857;
wire n_39_858;
wire n_39_859;
wire n_39_860;
wire n_39_861;
wire n_39_862;
wire \c1[28][31] ;
wire \c1[28][30] ;
wire \c1[28][29] ;
wire \c1[28][28] ;
wire \c1[28][27] ;
wire \c1[28][26] ;
wire \c1[28][25] ;
wire \c1[28][24] ;
wire \c1[28][23] ;
wire \c1[28][22] ;
wire \c1[28][21] ;
wire \c1[28][20] ;
wire \c1[28][19] ;
wire \c1[28][18] ;
wire \c1[28][17] ;
wire \c1[28][16] ;
wire \c1[28][15] ;
wire \c1[28][14] ;
wire \c1[28][13] ;
wire \c1[28][12] ;
wire \c1[28][11] ;
wire \c1[28][10] ;
wire \c1[28][9] ;
wire \c1[28][8] ;
wire \c1[28][7] ;
wire \c1[28][6] ;
wire \c1[28][5] ;
wire \c1[28][4] ;
wire \c1[28][3] ;
wire \c1[28][2] ;
wire \c1[28][1] ;
wire \c1[28][0] ;
wire n_39_864;
wire n_39_865;
wire n_39_866;
wire n_39_867;
wire n_39_31;
wire n_39_63;
wire n_39_95;
wire n_39_127;
wire n_39_159;
wire n_39_191;
wire n_39_223;
wire n_39_255;
wire n_39_287;
wire n_39_319;
wire n_39_351;
wire n_39_383;
wire n_39_415;
wire n_39_447;
wire n_39_479;
wire n_39_511;
wire n_39_543;
wire n_39_575;
wire n_39_607;
wire n_39_639;
wire n_39_671;
wire n_39_703;
wire n_39_735;
wire n_39_767;
wire n_39_799;
wire n_39_831;
wire n_39_863;
wire \c1[29][31] ;
wire \c1[29][30] ;
wire \c1[29][29] ;
wire \c1[29][28] ;
wire \c1[29][27] ;
wire \c1[29][26] ;
wire \c1[29][25] ;
wire \c1[29][24] ;
wire \c1[29][23] ;
wire \c1[29][22] ;
wire \c1[29][21] ;
wire \c1[29][20] ;
wire \c1[29][19] ;
wire \c1[29][18] ;
wire \c1[29][17] ;
wire \c1[29][16] ;
wire \c1[29][15] ;
wire \c1[29][14] ;
wire \c1[29][13] ;
wire \c1[29][12] ;
wire \c1[29][11] ;
wire \c1[29][10] ;
wire \c1[29][9] ;
wire \c1[29][8] ;
wire \c1[29][7] ;
wire \c1[29][6] ;
wire \c1[29][5] ;
wire \c1[29][4] ;
wire \c1[29][3] ;
wire \c1[29][2] ;
wire \c1[29][1] ;
wire \c1[29][0] ;
wire \s1[29][31] ;
wire \s1[29][30] ;
wire \s1[29][29] ;
wire \s1[29][28] ;
wire \s1[29][27] ;
wire \s1[29][26] ;
wire \s1[29][25] ;
wire \s1[29][24] ;
wire \s1[29][23] ;
wire \s1[29][22] ;
wire \s1[29][21] ;
wire \s1[29][20] ;
wire \s1[29][19] ;
wire \s1[29][18] ;
wire \s1[29][17] ;
wire \s1[29][16] ;
wire \s1[29][15] ;
wire \s1[29][14] ;
wire \s1[29][13] ;
wire \s1[29][12] ;
wire \s1[29][11] ;
wire \s1[29][10] ;
wire \s1[29][9] ;
wire \s1[29][8] ;
wire \s1[29][7] ;
wire \s1[29][6] ;
wire \s1[29][5] ;
wire \s1[29][4] ;
wire \s1[29][3] ;
wire \s1[29][2] ;
wire \s1[29][1] ;
wire \s1[29][0] ;
wire n_4_0_1;
wire n_4_0_2;
wire \partial_reg[0][31] ;
wire \partial_reg[0][30] ;
wire \partial_reg[0][29] ;
wire \partial_reg[0][28] ;
wire \partial_reg[0][27] ;
wire \partial_reg[0][26] ;
wire \partial_reg[0][25] ;
wire \partial_reg[0][24] ;
wire \partial_reg[0][23] ;
wire \partial_reg[0][22] ;
wire \partial_reg[0][21] ;
wire \partial_reg[0][20] ;
wire \partial_reg[0][19] ;
wire \partial_reg[0][18] ;
wire \partial_reg[0][17] ;
wire \partial_reg[0][16] ;
wire \partial_reg[0][15] ;
wire \partial_reg[0][14] ;
wire \partial_reg[0][13] ;
wire \partial_reg[0][12] ;
wire \partial_reg[0][11] ;
wire \partial_reg[0][10] ;
wire \partial_reg[0][9] ;
wire \partial_reg[0][8] ;
wire \partial_reg[0][7] ;
wire \partial_reg[0][6] ;
wire \partial_reg[0][5] ;
wire \partial_reg[0][4] ;
wire \partial_reg[0][3] ;
wire \partial_reg[0][2] ;
wire \partial_reg[0][1] ;
wire n_4_0_3;
wire n_4_0_4;
wire n_4_0_5;
wire n_4_0_6;
wire n_4_0_7;
wire n_4_0_8;
wire n_4_0_9;
wire n_4_0_10;
wire n_4_0_11;
wire n_4_0_12;
wire n_4_0_13;
wire n_4_0_14;
wire n_4_0_15;
wire n_4_0_16;
wire n_4_0_17;
wire n_4_0_18;
wire n_4_0_19;
wire n_4_0_20;
wire n_4_0_21;
wire n_4_0_22;
wire n_4_0_23;
wire n_4_0_24;
wire n_4_0_25;
wire n_4_0_26;
wire n_4_0_27;
wire n_4_0_28;
wire n_4_0_29;
wire \partial_reg[1][31] ;
wire \partial_reg[1][30] ;
wire \partial_reg[1][29] ;
wire \partial_reg[1][28] ;
wire \partial_reg[1][27] ;
wire \partial_reg[1][26] ;
wire \partial_reg[1][25] ;
wire \partial_reg[1][24] ;
wire \partial_reg[1][23] ;
wire \partial_reg[1][22] ;
wire \partial_reg[1][21] ;
wire \partial_reg[1][20] ;
wire \partial_reg[1][19] ;
wire \partial_reg[1][18] ;
wire \partial_reg[1][17] ;
wire \partial_reg[1][16] ;
wire \partial_reg[1][15] ;
wire \partial_reg[1][14] ;
wire \partial_reg[1][13] ;
wire \partial_reg[1][12] ;
wire \partial_reg[1][11] ;
wire \partial_reg[1][10] ;
wire \partial_reg[1][9] ;
wire \partial_reg[1][8] ;
wire \partial_reg[1][7] ;
wire \partial_reg[1][6] ;
wire \partial_reg[1][5] ;
wire \partial_reg[1][4] ;
wire \partial_reg[1][3] ;
wire \partial_reg[1][2] ;
wire \partial_reg[1][1] ;
wire \partial_reg[1][0] ;
wire \partial_reg[2][31] ;
wire \partial_reg[2][30] ;
wire \partial_reg[2][29] ;
wire \partial_reg[2][28] ;
wire \partial_reg[2][27] ;
wire \partial_reg[2][26] ;
wire \partial_reg[2][25] ;
wire \partial_reg[2][24] ;
wire \partial_reg[2][23] ;
wire \partial_reg[2][22] ;
wire \partial_reg[2][21] ;
wire \partial_reg[2][20] ;
wire \partial_reg[2][19] ;
wire \partial_reg[2][18] ;
wire \partial_reg[2][17] ;
wire \partial_reg[2][16] ;
wire \partial_reg[2][15] ;
wire \partial_reg[2][14] ;
wire \partial_reg[2][13] ;
wire \partial_reg[2][12] ;
wire \partial_reg[2][11] ;
wire \partial_reg[2][10] ;
wire \partial_reg[2][9] ;
wire \partial_reg[2][8] ;
wire \partial_reg[2][7] ;
wire \partial_reg[2][6] ;
wire \partial_reg[2][5] ;
wire \partial_reg[2][4] ;
wire \partial_reg[2][3] ;
wire \partial_reg[2][2] ;
wire \partial_reg[2][1] ;
wire \partial_reg[2][0] ;
wire n_4_0_35;
wire \partial_reg[3][31] ;
wire \partial_reg[3][30] ;
wire \partial_reg[3][29] ;
wire \partial_reg[3][28] ;
wire \partial_reg[3][27] ;
wire \partial_reg[3][26] ;
wire \partial_reg[3][25] ;
wire \partial_reg[3][24] ;
wire \partial_reg[3][23] ;
wire \partial_reg[3][22] ;
wire \partial_reg[3][21] ;
wire \partial_reg[3][20] ;
wire \partial_reg[3][19] ;
wire \partial_reg[3][18] ;
wire \partial_reg[3][17] ;
wire \partial_reg[3][16] ;
wire \partial_reg[3][15] ;
wire \partial_reg[3][14] ;
wire \partial_reg[3][13] ;
wire \partial_reg[3][12] ;
wire \partial_reg[3][11] ;
wire \partial_reg[3][10] ;
wire \partial_reg[3][9] ;
wire \partial_reg[3][8] ;
wire \partial_reg[3][7] ;
wire \partial_reg[3][6] ;
wire \partial_reg[3][5] ;
wire \partial_reg[3][4] ;
wire \partial_reg[3][3] ;
wire \partial_reg[3][2] ;
wire \partial_reg[3][1] ;
wire \partial_reg[3][0] ;
wire n_4_0_36;
wire \partial_reg[4][31] ;
wire \partial_reg[4][30] ;
wire \partial_reg[4][29] ;
wire \partial_reg[4][28] ;
wire \partial_reg[4][27] ;
wire \partial_reg[4][26] ;
wire \partial_reg[4][25] ;
wire \partial_reg[4][24] ;
wire \partial_reg[4][23] ;
wire \partial_reg[4][22] ;
wire \partial_reg[4][21] ;
wire \partial_reg[4][20] ;
wire \partial_reg[4][19] ;
wire \partial_reg[4][18] ;
wire \partial_reg[4][17] ;
wire \partial_reg[4][16] ;
wire \partial_reg[4][15] ;
wire \partial_reg[4][14] ;
wire \partial_reg[4][13] ;
wire \partial_reg[4][12] ;
wire \partial_reg[4][11] ;
wire \partial_reg[4][10] ;
wire \partial_reg[4][9] ;
wire \partial_reg[4][8] ;
wire \partial_reg[4][7] ;
wire \partial_reg[4][6] ;
wire \partial_reg[4][5] ;
wire \partial_reg[4][4] ;
wire \partial_reg[4][3] ;
wire \partial_reg[4][2] ;
wire \partial_reg[4][1] ;
wire \partial_reg[4][0] ;
wire n_4_0_37;
wire \partial_reg[5][31] ;
wire \partial_reg[5][30] ;
wire \partial_reg[5][29] ;
wire \partial_reg[5][28] ;
wire \partial_reg[5][27] ;
wire \partial_reg[5][26] ;
wire \partial_reg[5][25] ;
wire \partial_reg[5][24] ;
wire \partial_reg[5][23] ;
wire \partial_reg[5][22] ;
wire \partial_reg[5][21] ;
wire \partial_reg[5][20] ;
wire \partial_reg[5][19] ;
wire \partial_reg[5][18] ;
wire \partial_reg[5][17] ;
wire \partial_reg[5][16] ;
wire \partial_reg[5][15] ;
wire \partial_reg[5][14] ;
wire \partial_reg[5][13] ;
wire \partial_reg[5][12] ;
wire \partial_reg[5][11] ;
wire \partial_reg[5][10] ;
wire \partial_reg[5][9] ;
wire \partial_reg[5][8] ;
wire \partial_reg[5][7] ;
wire \partial_reg[5][6] ;
wire \partial_reg[5][5] ;
wire \partial_reg[5][4] ;
wire \partial_reg[5][3] ;
wire \partial_reg[5][2] ;
wire \partial_reg[5][1] ;
wire \partial_reg[5][0] ;
wire n_4_0_38;
wire \partial_reg[6][31] ;
wire \partial_reg[6][30] ;
wire \partial_reg[6][29] ;
wire \partial_reg[6][28] ;
wire \partial_reg[6][27] ;
wire \partial_reg[6][26] ;
wire \partial_reg[6][25] ;
wire \partial_reg[6][24] ;
wire \partial_reg[6][23] ;
wire \partial_reg[6][22] ;
wire \partial_reg[6][21] ;
wire \partial_reg[6][20] ;
wire \partial_reg[6][19] ;
wire \partial_reg[6][18] ;
wire \partial_reg[6][17] ;
wire \partial_reg[6][16] ;
wire \partial_reg[6][15] ;
wire \partial_reg[6][14] ;
wire \partial_reg[6][13] ;
wire \partial_reg[6][12] ;
wire \partial_reg[6][11] ;
wire \partial_reg[6][10] ;
wire \partial_reg[6][9] ;
wire \partial_reg[6][8] ;
wire \partial_reg[6][7] ;
wire \partial_reg[6][6] ;
wire \partial_reg[6][5] ;
wire \partial_reg[6][4] ;
wire \partial_reg[6][3] ;
wire \partial_reg[6][2] ;
wire \partial_reg[6][1] ;
wire \partial_reg[6][0] ;
wire n_4_0_39;
wire \partial_reg[7][31] ;
wire \partial_reg[7][30] ;
wire \partial_reg[7][29] ;
wire \partial_reg[7][28] ;
wire \partial_reg[7][27] ;
wire \partial_reg[7][26] ;
wire \partial_reg[7][25] ;
wire \partial_reg[7][24] ;
wire \partial_reg[7][23] ;
wire \partial_reg[7][22] ;
wire \partial_reg[7][21] ;
wire \partial_reg[7][20] ;
wire \partial_reg[7][19] ;
wire \partial_reg[7][18] ;
wire \partial_reg[7][17] ;
wire \partial_reg[7][16] ;
wire \partial_reg[7][15] ;
wire \partial_reg[7][14] ;
wire \partial_reg[7][13] ;
wire \partial_reg[7][12] ;
wire \partial_reg[7][11] ;
wire \partial_reg[7][10] ;
wire \partial_reg[7][9] ;
wire \partial_reg[7][8] ;
wire \partial_reg[7][7] ;
wire \partial_reg[7][6] ;
wire \partial_reg[7][5] ;
wire \partial_reg[7][4] ;
wire \partial_reg[7][3] ;
wire \partial_reg[7][2] ;
wire \partial_reg[7][1] ;
wire \partial_reg[7][0] ;
wire n_4_0_40;
wire \partial_reg[8][31] ;
wire \partial_reg[8][30] ;
wire \partial_reg[8][29] ;
wire \partial_reg[8][28] ;
wire \partial_reg[8][27] ;
wire \partial_reg[8][26] ;
wire \partial_reg[8][25] ;
wire \partial_reg[8][24] ;
wire \partial_reg[8][23] ;
wire \partial_reg[8][22] ;
wire \partial_reg[8][21] ;
wire \partial_reg[8][20] ;
wire \partial_reg[8][19] ;
wire \partial_reg[8][18] ;
wire \partial_reg[8][17] ;
wire \partial_reg[8][16] ;
wire \partial_reg[8][15] ;
wire \partial_reg[8][14] ;
wire \partial_reg[8][13] ;
wire \partial_reg[8][12] ;
wire \partial_reg[8][11] ;
wire \partial_reg[8][10] ;
wire \partial_reg[8][9] ;
wire \partial_reg[8][8] ;
wire \partial_reg[8][7] ;
wire \partial_reg[8][6] ;
wire \partial_reg[8][5] ;
wire \partial_reg[8][4] ;
wire \partial_reg[8][3] ;
wire \partial_reg[8][2] ;
wire \partial_reg[8][1] ;
wire \partial_reg[8][0] ;
wire n_4_0_41;
wire \partial_reg[9][31] ;
wire \partial_reg[9][30] ;
wire \partial_reg[9][29] ;
wire \partial_reg[9][28] ;
wire \partial_reg[9][27] ;
wire \partial_reg[9][26] ;
wire \partial_reg[9][25] ;
wire \partial_reg[9][24] ;
wire \partial_reg[9][23] ;
wire \partial_reg[9][22] ;
wire \partial_reg[9][21] ;
wire \partial_reg[9][20] ;
wire \partial_reg[9][19] ;
wire \partial_reg[9][18] ;
wire \partial_reg[9][17] ;
wire \partial_reg[9][16] ;
wire \partial_reg[9][15] ;
wire \partial_reg[9][14] ;
wire \partial_reg[9][13] ;
wire \partial_reg[9][12] ;
wire \partial_reg[9][11] ;
wire \partial_reg[9][10] ;
wire \partial_reg[9][9] ;
wire \partial_reg[9][8] ;
wire \partial_reg[9][7] ;
wire \partial_reg[9][6] ;
wire \partial_reg[9][5] ;
wire \partial_reg[9][4] ;
wire \partial_reg[9][3] ;
wire \partial_reg[9][2] ;
wire \partial_reg[9][1] ;
wire \partial_reg[9][0] ;
wire n_4_0_42;
wire \partial_reg[10][31] ;
wire \partial_reg[10][30] ;
wire \partial_reg[10][29] ;
wire \partial_reg[10][28] ;
wire \partial_reg[10][27] ;
wire \partial_reg[10][26] ;
wire \partial_reg[10][25] ;
wire \partial_reg[10][24] ;
wire \partial_reg[10][23] ;
wire \partial_reg[10][22] ;
wire \partial_reg[10][21] ;
wire \partial_reg[10][20] ;
wire \partial_reg[10][19] ;
wire \partial_reg[10][18] ;
wire \partial_reg[10][17] ;
wire \partial_reg[10][16] ;
wire \partial_reg[10][15] ;
wire \partial_reg[10][14] ;
wire \partial_reg[10][13] ;
wire \partial_reg[10][12] ;
wire \partial_reg[10][11] ;
wire \partial_reg[10][10] ;
wire \partial_reg[10][9] ;
wire \partial_reg[10][8] ;
wire \partial_reg[10][7] ;
wire \partial_reg[10][6] ;
wire \partial_reg[10][5] ;
wire \partial_reg[10][4] ;
wire \partial_reg[10][3] ;
wire \partial_reg[10][2] ;
wire \partial_reg[10][1] ;
wire \partial_reg[10][0] ;
wire n_4_0_43;
wire \partial_reg[11][31] ;
wire \partial_reg[11][30] ;
wire \partial_reg[11][29] ;
wire \partial_reg[11][28] ;
wire \partial_reg[11][27] ;
wire \partial_reg[11][26] ;
wire \partial_reg[11][25] ;
wire \partial_reg[11][24] ;
wire \partial_reg[11][23] ;
wire \partial_reg[11][22] ;
wire \partial_reg[11][21] ;
wire \partial_reg[11][20] ;
wire \partial_reg[11][19] ;
wire \partial_reg[11][18] ;
wire \partial_reg[11][17] ;
wire \partial_reg[11][16] ;
wire \partial_reg[11][15] ;
wire \partial_reg[11][14] ;
wire \partial_reg[11][13] ;
wire \partial_reg[11][12] ;
wire \partial_reg[11][11] ;
wire \partial_reg[11][10] ;
wire \partial_reg[11][9] ;
wire \partial_reg[11][8] ;
wire \partial_reg[11][7] ;
wire \partial_reg[11][6] ;
wire \partial_reg[11][5] ;
wire \partial_reg[11][4] ;
wire \partial_reg[11][3] ;
wire \partial_reg[11][2] ;
wire \partial_reg[11][1] ;
wire \partial_reg[11][0] ;
wire n_4_0_44;
wire \partial_reg[12][31] ;
wire \partial_reg[12][30] ;
wire \partial_reg[12][29] ;
wire \partial_reg[12][28] ;
wire \partial_reg[12][27] ;
wire \partial_reg[12][26] ;
wire \partial_reg[12][25] ;
wire \partial_reg[12][24] ;
wire \partial_reg[12][23] ;
wire \partial_reg[12][22] ;
wire \partial_reg[12][21] ;
wire \partial_reg[12][20] ;
wire \partial_reg[12][19] ;
wire \partial_reg[12][18] ;
wire \partial_reg[12][17] ;
wire \partial_reg[12][16] ;
wire \partial_reg[12][15] ;
wire \partial_reg[12][14] ;
wire \partial_reg[12][13] ;
wire \partial_reg[12][12] ;
wire \partial_reg[12][11] ;
wire \partial_reg[12][10] ;
wire \partial_reg[12][9] ;
wire \partial_reg[12][8] ;
wire \partial_reg[12][7] ;
wire \partial_reg[12][6] ;
wire \partial_reg[12][5] ;
wire \partial_reg[12][4] ;
wire \partial_reg[12][3] ;
wire \partial_reg[12][2] ;
wire \partial_reg[12][1] ;
wire \partial_reg[12][0] ;
wire n_4_0_45;
wire \partial_reg[13][31] ;
wire \partial_reg[13][30] ;
wire \partial_reg[13][29] ;
wire \partial_reg[13][28] ;
wire \partial_reg[13][27] ;
wire \partial_reg[13][26] ;
wire \partial_reg[13][25] ;
wire \partial_reg[13][24] ;
wire \partial_reg[13][23] ;
wire \partial_reg[13][22] ;
wire \partial_reg[13][21] ;
wire \partial_reg[13][20] ;
wire \partial_reg[13][19] ;
wire \partial_reg[13][18] ;
wire \partial_reg[13][17] ;
wire \partial_reg[13][16] ;
wire \partial_reg[13][15] ;
wire \partial_reg[13][14] ;
wire \partial_reg[13][13] ;
wire \partial_reg[13][12] ;
wire \partial_reg[13][11] ;
wire \partial_reg[13][10] ;
wire \partial_reg[13][9] ;
wire \partial_reg[13][8] ;
wire \partial_reg[13][7] ;
wire \partial_reg[13][6] ;
wire \partial_reg[13][5] ;
wire \partial_reg[13][4] ;
wire \partial_reg[13][3] ;
wire \partial_reg[13][2] ;
wire \partial_reg[13][1] ;
wire \partial_reg[13][0] ;
wire n_4_0_46;
wire \partial_reg[14][31] ;
wire \partial_reg[14][30] ;
wire \partial_reg[14][29] ;
wire \partial_reg[14][28] ;
wire \partial_reg[14][27] ;
wire \partial_reg[14][26] ;
wire \partial_reg[14][25] ;
wire \partial_reg[14][24] ;
wire \partial_reg[14][23] ;
wire \partial_reg[14][22] ;
wire \partial_reg[14][21] ;
wire \partial_reg[14][20] ;
wire \partial_reg[14][19] ;
wire \partial_reg[14][18] ;
wire \partial_reg[14][17] ;
wire \partial_reg[14][16] ;
wire \partial_reg[14][15] ;
wire \partial_reg[14][14] ;
wire \partial_reg[14][13] ;
wire \partial_reg[14][12] ;
wire \partial_reg[14][11] ;
wire \partial_reg[14][10] ;
wire \partial_reg[14][9] ;
wire \partial_reg[14][8] ;
wire \partial_reg[14][7] ;
wire \partial_reg[14][6] ;
wire \partial_reg[14][5] ;
wire \partial_reg[14][4] ;
wire \partial_reg[14][3] ;
wire \partial_reg[14][2] ;
wire \partial_reg[14][1] ;
wire \partial_reg[14][0] ;
wire n_4_0_47;
wire \partial_reg[15][31] ;
wire \partial_reg[15][30] ;
wire \partial_reg[15][29] ;
wire \partial_reg[15][28] ;
wire \partial_reg[15][27] ;
wire \partial_reg[15][26] ;
wire \partial_reg[15][25] ;
wire \partial_reg[15][24] ;
wire \partial_reg[15][23] ;
wire \partial_reg[15][22] ;
wire \partial_reg[15][21] ;
wire \partial_reg[15][20] ;
wire \partial_reg[15][19] ;
wire \partial_reg[15][18] ;
wire \partial_reg[15][17] ;
wire \partial_reg[15][16] ;
wire \partial_reg[15][15] ;
wire \partial_reg[15][14] ;
wire \partial_reg[15][13] ;
wire \partial_reg[15][12] ;
wire \partial_reg[15][11] ;
wire \partial_reg[15][10] ;
wire \partial_reg[15][9] ;
wire \partial_reg[15][8] ;
wire \partial_reg[15][7] ;
wire \partial_reg[15][6] ;
wire \partial_reg[15][5] ;
wire \partial_reg[15][4] ;
wire \partial_reg[15][3] ;
wire \partial_reg[15][2] ;
wire \partial_reg[15][1] ;
wire \partial_reg[15][0] ;
wire n_4_0_48;
wire \partial_reg[16][31] ;
wire \partial_reg[16][30] ;
wire \partial_reg[16][29] ;
wire \partial_reg[16][28] ;
wire \partial_reg[16][27] ;
wire \partial_reg[16][26] ;
wire \partial_reg[16][25] ;
wire \partial_reg[16][24] ;
wire \partial_reg[16][23] ;
wire \partial_reg[16][22] ;
wire \partial_reg[16][21] ;
wire \partial_reg[16][20] ;
wire \partial_reg[16][19] ;
wire \partial_reg[16][18] ;
wire \partial_reg[16][17] ;
wire \partial_reg[16][16] ;
wire \partial_reg[16][15] ;
wire \partial_reg[16][14] ;
wire \partial_reg[16][13] ;
wire \partial_reg[16][12] ;
wire \partial_reg[16][11] ;
wire \partial_reg[16][10] ;
wire \partial_reg[16][9] ;
wire \partial_reg[16][8] ;
wire \partial_reg[16][7] ;
wire \partial_reg[16][6] ;
wire \partial_reg[16][5] ;
wire \partial_reg[16][4] ;
wire \partial_reg[16][3] ;
wire \partial_reg[16][2] ;
wire \partial_reg[16][1] ;
wire \partial_reg[16][0] ;
wire n_4_0_49;
wire \partial_reg[17][31] ;
wire \partial_reg[17][30] ;
wire \partial_reg[17][29] ;
wire \partial_reg[17][28] ;
wire \partial_reg[17][27] ;
wire \partial_reg[17][26] ;
wire \partial_reg[17][25] ;
wire \partial_reg[17][24] ;
wire \partial_reg[17][23] ;
wire \partial_reg[17][22] ;
wire \partial_reg[17][21] ;
wire \partial_reg[17][20] ;
wire \partial_reg[17][19] ;
wire \partial_reg[17][18] ;
wire \partial_reg[17][17] ;
wire \partial_reg[17][16] ;
wire \partial_reg[17][15] ;
wire \partial_reg[17][14] ;
wire \partial_reg[17][13] ;
wire \partial_reg[17][12] ;
wire \partial_reg[17][11] ;
wire \partial_reg[17][10] ;
wire \partial_reg[17][9] ;
wire \partial_reg[17][8] ;
wire \partial_reg[17][7] ;
wire \partial_reg[17][6] ;
wire \partial_reg[17][5] ;
wire \partial_reg[17][4] ;
wire \partial_reg[17][3] ;
wire \partial_reg[17][2] ;
wire \partial_reg[17][1] ;
wire \partial_reg[17][0] ;
wire n_4_0_50;
wire \partial_reg[18][31] ;
wire \partial_reg[18][30] ;
wire \partial_reg[18][29] ;
wire \partial_reg[18][28] ;
wire \partial_reg[18][27] ;
wire \partial_reg[18][26] ;
wire \partial_reg[18][25] ;
wire \partial_reg[18][24] ;
wire \partial_reg[18][23] ;
wire \partial_reg[18][22] ;
wire \partial_reg[18][21] ;
wire \partial_reg[18][20] ;
wire \partial_reg[18][19] ;
wire \partial_reg[18][18] ;
wire \partial_reg[18][17] ;
wire \partial_reg[18][16] ;
wire \partial_reg[18][15] ;
wire \partial_reg[18][14] ;
wire \partial_reg[18][13] ;
wire \partial_reg[18][12] ;
wire \partial_reg[18][11] ;
wire \partial_reg[18][10] ;
wire \partial_reg[18][9] ;
wire \partial_reg[18][8] ;
wire \partial_reg[18][7] ;
wire \partial_reg[18][6] ;
wire \partial_reg[18][5] ;
wire \partial_reg[18][4] ;
wire \partial_reg[18][3] ;
wire \partial_reg[18][2] ;
wire \partial_reg[18][1] ;
wire \partial_reg[18][0] ;
wire n_4_0_51;
wire \partial_reg[19][31] ;
wire \partial_reg[19][30] ;
wire \partial_reg[19][29] ;
wire \partial_reg[19][28] ;
wire \partial_reg[19][27] ;
wire \partial_reg[19][26] ;
wire \partial_reg[19][25] ;
wire \partial_reg[19][24] ;
wire \partial_reg[19][23] ;
wire \partial_reg[19][22] ;
wire \partial_reg[19][21] ;
wire \partial_reg[19][20] ;
wire \partial_reg[19][19] ;
wire \partial_reg[19][18] ;
wire \partial_reg[19][17] ;
wire \partial_reg[19][16] ;
wire \partial_reg[19][15] ;
wire \partial_reg[19][14] ;
wire \partial_reg[19][13] ;
wire \partial_reg[19][12] ;
wire \partial_reg[19][11] ;
wire \partial_reg[19][10] ;
wire \partial_reg[19][9] ;
wire \partial_reg[19][8] ;
wire \partial_reg[19][7] ;
wire \partial_reg[19][6] ;
wire \partial_reg[19][5] ;
wire \partial_reg[19][4] ;
wire \partial_reg[19][3] ;
wire \partial_reg[19][2] ;
wire \partial_reg[19][1] ;
wire \partial_reg[19][0] ;
wire n_4_0_52;
wire \partial_reg[20][31] ;
wire \partial_reg[20][30] ;
wire \partial_reg[20][29] ;
wire \partial_reg[20][28] ;
wire \partial_reg[20][27] ;
wire \partial_reg[20][26] ;
wire \partial_reg[20][25] ;
wire \partial_reg[20][24] ;
wire \partial_reg[20][23] ;
wire \partial_reg[20][22] ;
wire \partial_reg[20][21] ;
wire \partial_reg[20][20] ;
wire \partial_reg[20][19] ;
wire \partial_reg[20][18] ;
wire \partial_reg[20][17] ;
wire \partial_reg[20][16] ;
wire \partial_reg[20][15] ;
wire \partial_reg[20][14] ;
wire \partial_reg[20][13] ;
wire \partial_reg[20][12] ;
wire \partial_reg[20][11] ;
wire \partial_reg[20][10] ;
wire \partial_reg[20][9] ;
wire \partial_reg[20][8] ;
wire \partial_reg[20][7] ;
wire \partial_reg[20][6] ;
wire \partial_reg[20][5] ;
wire \partial_reg[20][4] ;
wire \partial_reg[20][3] ;
wire \partial_reg[20][2] ;
wire \partial_reg[20][1] ;
wire \partial_reg[20][0] ;
wire n_4_0_53;
wire \partial_reg[21][31] ;
wire \partial_reg[21][30] ;
wire \partial_reg[21][29] ;
wire \partial_reg[21][28] ;
wire \partial_reg[21][27] ;
wire \partial_reg[21][26] ;
wire \partial_reg[21][25] ;
wire \partial_reg[21][24] ;
wire \partial_reg[21][23] ;
wire \partial_reg[21][22] ;
wire \partial_reg[21][21] ;
wire \partial_reg[21][20] ;
wire \partial_reg[21][19] ;
wire \partial_reg[21][18] ;
wire \partial_reg[21][17] ;
wire \partial_reg[21][16] ;
wire \partial_reg[21][15] ;
wire \partial_reg[21][14] ;
wire \partial_reg[21][13] ;
wire \partial_reg[21][12] ;
wire \partial_reg[21][11] ;
wire \partial_reg[21][10] ;
wire \partial_reg[21][9] ;
wire \partial_reg[21][8] ;
wire \partial_reg[21][7] ;
wire \partial_reg[21][6] ;
wire \partial_reg[21][5] ;
wire \partial_reg[21][4] ;
wire \partial_reg[21][3] ;
wire \partial_reg[21][2] ;
wire \partial_reg[21][1] ;
wire \partial_reg[21][0] ;
wire n_4_0_54;
wire \partial_reg[22][31] ;
wire \partial_reg[22][30] ;
wire \partial_reg[22][29] ;
wire \partial_reg[22][28] ;
wire \partial_reg[22][27] ;
wire \partial_reg[22][26] ;
wire \partial_reg[22][25] ;
wire \partial_reg[22][24] ;
wire \partial_reg[22][23] ;
wire \partial_reg[22][22] ;
wire \partial_reg[22][21] ;
wire \partial_reg[22][20] ;
wire \partial_reg[22][19] ;
wire \partial_reg[22][18] ;
wire \partial_reg[22][17] ;
wire \partial_reg[22][16] ;
wire \partial_reg[22][15] ;
wire \partial_reg[22][14] ;
wire \partial_reg[22][13] ;
wire \partial_reg[22][12] ;
wire \partial_reg[22][11] ;
wire \partial_reg[22][10] ;
wire \partial_reg[22][9] ;
wire \partial_reg[22][8] ;
wire \partial_reg[22][7] ;
wire \partial_reg[22][6] ;
wire \partial_reg[22][5] ;
wire \partial_reg[22][4] ;
wire \partial_reg[22][3] ;
wire \partial_reg[22][2] ;
wire \partial_reg[22][1] ;
wire \partial_reg[22][0] ;
wire n_4_0_55;
wire \partial_reg[23][31] ;
wire \partial_reg[23][30] ;
wire \partial_reg[23][29] ;
wire \partial_reg[23][28] ;
wire \partial_reg[23][27] ;
wire \partial_reg[23][26] ;
wire \partial_reg[23][25] ;
wire \partial_reg[23][24] ;
wire \partial_reg[23][23] ;
wire \partial_reg[23][22] ;
wire \partial_reg[23][21] ;
wire \partial_reg[23][20] ;
wire \partial_reg[23][19] ;
wire \partial_reg[23][18] ;
wire \partial_reg[23][17] ;
wire \partial_reg[23][16] ;
wire \partial_reg[23][15] ;
wire \partial_reg[23][14] ;
wire \partial_reg[23][13] ;
wire \partial_reg[23][12] ;
wire \partial_reg[23][11] ;
wire \partial_reg[23][10] ;
wire \partial_reg[23][9] ;
wire \partial_reg[23][8] ;
wire \partial_reg[23][7] ;
wire \partial_reg[23][6] ;
wire \partial_reg[23][5] ;
wire \partial_reg[23][4] ;
wire \partial_reg[23][3] ;
wire \partial_reg[23][2] ;
wire \partial_reg[23][1] ;
wire \partial_reg[23][0] ;
wire n_4_0_56;
wire \partial_reg[24][31] ;
wire \partial_reg[24][30] ;
wire \partial_reg[24][29] ;
wire \partial_reg[24][28] ;
wire \partial_reg[24][27] ;
wire \partial_reg[24][26] ;
wire \partial_reg[24][25] ;
wire \partial_reg[24][24] ;
wire \partial_reg[24][23] ;
wire \partial_reg[24][22] ;
wire \partial_reg[24][21] ;
wire \partial_reg[24][20] ;
wire \partial_reg[24][19] ;
wire \partial_reg[24][18] ;
wire \partial_reg[24][17] ;
wire \partial_reg[24][16] ;
wire \partial_reg[24][15] ;
wire \partial_reg[24][14] ;
wire \partial_reg[24][13] ;
wire \partial_reg[24][12] ;
wire \partial_reg[24][11] ;
wire \partial_reg[24][10] ;
wire \partial_reg[24][9] ;
wire \partial_reg[24][8] ;
wire \partial_reg[24][7] ;
wire \partial_reg[24][6] ;
wire \partial_reg[24][5] ;
wire \partial_reg[24][4] ;
wire \partial_reg[24][3] ;
wire \partial_reg[24][2] ;
wire \partial_reg[24][1] ;
wire \partial_reg[24][0] ;
wire n_4_0_57;
wire \partial_reg[25][31] ;
wire \partial_reg[25][30] ;
wire \partial_reg[25][29] ;
wire \partial_reg[25][28] ;
wire \partial_reg[25][27] ;
wire \partial_reg[25][26] ;
wire \partial_reg[25][25] ;
wire \partial_reg[25][24] ;
wire \partial_reg[25][23] ;
wire \partial_reg[25][22] ;
wire \partial_reg[25][21] ;
wire \partial_reg[25][20] ;
wire \partial_reg[25][19] ;
wire \partial_reg[25][18] ;
wire \partial_reg[25][17] ;
wire \partial_reg[25][16] ;
wire \partial_reg[25][15] ;
wire \partial_reg[25][14] ;
wire \partial_reg[25][13] ;
wire \partial_reg[25][12] ;
wire \partial_reg[25][11] ;
wire \partial_reg[25][10] ;
wire \partial_reg[25][9] ;
wire \partial_reg[25][8] ;
wire \partial_reg[25][7] ;
wire \partial_reg[25][6] ;
wire \partial_reg[25][5] ;
wire \partial_reg[25][4] ;
wire \partial_reg[25][3] ;
wire \partial_reg[25][2] ;
wire \partial_reg[25][1] ;
wire \partial_reg[25][0] ;
wire n_4_0_58;
wire \partial_reg[26][31] ;
wire \partial_reg[26][30] ;
wire \partial_reg[26][29] ;
wire \partial_reg[26][28] ;
wire \partial_reg[26][27] ;
wire \partial_reg[26][26] ;
wire \partial_reg[26][25] ;
wire \partial_reg[26][24] ;
wire \partial_reg[26][23] ;
wire \partial_reg[26][22] ;
wire \partial_reg[26][21] ;
wire \partial_reg[26][20] ;
wire \partial_reg[26][19] ;
wire \partial_reg[26][18] ;
wire \partial_reg[26][17] ;
wire \partial_reg[26][16] ;
wire \partial_reg[26][15] ;
wire \partial_reg[26][14] ;
wire \partial_reg[26][13] ;
wire \partial_reg[26][12] ;
wire \partial_reg[26][11] ;
wire \partial_reg[26][10] ;
wire \partial_reg[26][9] ;
wire \partial_reg[26][8] ;
wire \partial_reg[26][7] ;
wire \partial_reg[26][6] ;
wire \partial_reg[26][5] ;
wire \partial_reg[26][4] ;
wire \partial_reg[26][3] ;
wire \partial_reg[26][2] ;
wire \partial_reg[26][1] ;
wire \partial_reg[26][0] ;
wire n_4_0_59;
wire \partial_reg[27][31] ;
wire \partial_reg[27][30] ;
wire \partial_reg[27][29] ;
wire \partial_reg[27][28] ;
wire \partial_reg[27][27] ;
wire \partial_reg[27][26] ;
wire \partial_reg[27][25] ;
wire \partial_reg[27][24] ;
wire \partial_reg[27][23] ;
wire \partial_reg[27][22] ;
wire \partial_reg[27][21] ;
wire \partial_reg[27][20] ;
wire \partial_reg[27][19] ;
wire \partial_reg[27][18] ;
wire \partial_reg[27][17] ;
wire \partial_reg[27][16] ;
wire \partial_reg[27][15] ;
wire \partial_reg[27][14] ;
wire \partial_reg[27][13] ;
wire \partial_reg[27][12] ;
wire \partial_reg[27][11] ;
wire \partial_reg[27][10] ;
wire \partial_reg[27][9] ;
wire \partial_reg[27][8] ;
wire \partial_reg[27][7] ;
wire \partial_reg[27][6] ;
wire \partial_reg[27][5] ;
wire \partial_reg[27][4] ;
wire \partial_reg[27][3] ;
wire \partial_reg[27][2] ;
wire \partial_reg[27][1] ;
wire \partial_reg[27][0] ;
wire n_4_0_60;
wire \partial_reg[28][31] ;
wire \partial_reg[28][30] ;
wire \partial_reg[28][29] ;
wire \partial_reg[28][28] ;
wire \partial_reg[28][27] ;
wire \partial_reg[28][26] ;
wire \partial_reg[28][25] ;
wire \partial_reg[28][24] ;
wire \partial_reg[28][23] ;
wire \partial_reg[28][22] ;
wire \partial_reg[28][21] ;
wire \partial_reg[28][20] ;
wire \partial_reg[28][19] ;
wire \partial_reg[28][18] ;
wire \partial_reg[28][17] ;
wire \partial_reg[28][16] ;
wire \partial_reg[28][15] ;
wire \partial_reg[28][14] ;
wire \partial_reg[28][13] ;
wire \partial_reg[28][12] ;
wire \partial_reg[28][11] ;
wire \partial_reg[28][10] ;
wire \partial_reg[28][9] ;
wire \partial_reg[28][8] ;
wire \partial_reg[28][7] ;
wire \partial_reg[28][6] ;
wire \partial_reg[28][5] ;
wire \partial_reg[28][4] ;
wire \partial_reg[28][3] ;
wire \partial_reg[28][2] ;
wire \partial_reg[28][1] ;
wire \partial_reg[28][0] ;
wire n_4_0_61;
wire \partial_reg[29][31] ;
wire \partial_reg[29][30] ;
wire \partial_reg[29][29] ;
wire \partial_reg[29][28] ;
wire \partial_reg[29][27] ;
wire \partial_reg[29][26] ;
wire \partial_reg[29][25] ;
wire \partial_reg[29][24] ;
wire \partial_reg[29][23] ;
wire \partial_reg[29][22] ;
wire \partial_reg[29][21] ;
wire \partial_reg[29][20] ;
wire \partial_reg[29][19] ;
wire \partial_reg[29][18] ;
wire \partial_reg[29][17] ;
wire \partial_reg[29][16] ;
wire \partial_reg[29][15] ;
wire \partial_reg[29][14] ;
wire \partial_reg[29][13] ;
wire \partial_reg[29][12] ;
wire \partial_reg[29][11] ;
wire \partial_reg[29][10] ;
wire \partial_reg[29][9] ;
wire \partial_reg[29][8] ;
wire \partial_reg[29][7] ;
wire \partial_reg[29][6] ;
wire \partial_reg[29][5] ;
wire \partial_reg[29][4] ;
wire \partial_reg[29][3] ;
wire \partial_reg[29][2] ;
wire \partial_reg[29][1] ;
wire \partial_reg[29][0] ;
wire n_4_0_62;
wire \partial_reg[30][31] ;
wire \partial_reg[30][30] ;
wire \partial_reg[30][29] ;
wire \partial_reg[30][28] ;
wire \partial_reg[30][27] ;
wire \partial_reg[30][26] ;
wire \partial_reg[30][25] ;
wire \partial_reg[30][24] ;
wire \partial_reg[30][23] ;
wire \partial_reg[30][22] ;
wire \partial_reg[30][21] ;
wire \partial_reg[30][20] ;
wire \partial_reg[30][19] ;
wire \partial_reg[30][18] ;
wire \partial_reg[30][17] ;
wire \partial_reg[30][16] ;
wire \partial_reg[30][15] ;
wire \partial_reg[30][14] ;
wire \partial_reg[30][13] ;
wire \partial_reg[30][12] ;
wire \partial_reg[30][11] ;
wire \partial_reg[30][10] ;
wire \partial_reg[30][9] ;
wire \partial_reg[30][8] ;
wire \partial_reg[30][7] ;
wire \partial_reg[30][6] ;
wire \partial_reg[30][5] ;
wire \partial_reg[30][4] ;
wire \partial_reg[30][3] ;
wire \partial_reg[30][2] ;
wire \partial_reg[30][1] ;
wire \partial_reg[30][0] ;
wire n_4_0_63;
wire \partial_reg[31][31] ;
wire \partial_reg[31][30] ;
wire \partial_reg[31][29] ;
wire \partial_reg[31][28] ;
wire \partial_reg[31][27] ;
wire \partial_reg[31][26] ;
wire \partial_reg[31][25] ;
wire \partial_reg[31][24] ;
wire \partial_reg[31][23] ;
wire \partial_reg[31][22] ;
wire \partial_reg[31][21] ;
wire \partial_reg[31][20] ;
wire \partial_reg[31][19] ;
wire \partial_reg[31][18] ;
wire \partial_reg[31][17] ;
wire \partial_reg[31][16] ;
wire \partial_reg[31][15] ;
wire \partial_reg[31][14] ;
wire \partial_reg[31][13] ;
wire \partial_reg[31][12] ;
wire \partial_reg[31][11] ;
wire \partial_reg[31][10] ;
wire \partial_reg[31][9] ;
wire \partial_reg[31][8] ;
wire \partial_reg[31][7] ;
wire \partial_reg[31][6] ;
wire \partial_reg[31][5] ;
wire \partial_reg[31][4] ;
wire \partial_reg[31][3] ;
wire \partial_reg[31][2] ;
wire \partial_reg[31][1] ;
wire \partial_reg[31][0] ;
wire n_4_0_34;
wire n_4_0_33;
wire n_4_0_32;
wire n_4_0_31;
wire n_4_0_30;
wire n_4_0_0;
wire n_4_0_64;
wire n_4_0_65;
wire \c1[0][31] ;
wire \c1[0][30] ;
wire \c1[0][29] ;
wire \c1[0][28] ;
wire \c1[0][27] ;
wire \c1[0][26] ;
wire \c1[0][25] ;
wire \c1[0][24] ;
wire \c1[0][23] ;
wire \c1[0][22] ;
wire \c1[0][21] ;
wire \c1[0][20] ;
wire \c1[0][19] ;
wire \c1[0][18] ;
wire \c1[0][17] ;
wire \c1[0][16] ;
wire \c1[0][15] ;
wire \c1[0][14] ;
wire \c1[0][13] ;
wire \c1[0][12] ;
wire \c1[0][11] ;
wire \c1[0][10] ;
wire \c1[0][9] ;
wire \c1[0][8] ;
wire \c1[0][7] ;
wire \c1[0][6] ;
wire \c1[0][5] ;
wire \c1[0][4] ;
wire \c1[0][3] ;
wire \c1[0][2] ;
wire \c1[0][1] ;
wire \c1[0][0] ;
wire \s1[0][31] ;
wire \s1[0][30] ;
wire \s1[0][29] ;
wire \s1[0][28] ;
wire \s1[0][27] ;
wire \s1[0][26] ;
wire \s1[0][25] ;
wire \s1[0][24] ;
wire \s1[0][23] ;
wire \s1[0][22] ;
wire \s1[0][21] ;
wire \s1[0][20] ;
wire \s1[0][19] ;
wire \s1[0][18] ;
wire \s1[0][17] ;
wire \s1[0][16] ;
wire \s1[0][15] ;
wire \s1[0][14] ;
wire \s1[0][13] ;
wire \s1[0][12] ;
wire \s1[0][11] ;
wire \s1[0][10] ;
wire \s1[0][9] ;
wire \s1[0][8] ;
wire \s1[0][7] ;
wire \s1[0][6] ;
wire \s1[0][5] ;
wire \s1[0][4] ;
wire \s1[0][3] ;
wire \s1[0][2] ;
wire \s1[0][1] ;
wire \s1[0][0] ;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire \op2[31] ;
wire \op2[30] ;
wire \op2[29] ;
wire \op2[28] ;
wire \op2[27] ;
wire \op2[26] ;
wire \op2[25] ;
wire \op2[24] ;
wire \op2[23] ;
wire \op2[22] ;
wire \op2[21] ;
wire \op2[20] ;
wire \op2[19] ;
wire \op2[18] ;
wire \op2[17] ;
wire \op2[16] ;
wire \op2[15] ;
wire \op2[14] ;
wire \op2[13] ;
wire \op2[12] ;
wire \op2[11] ;
wire \op2[10] ;
wire \op2[9] ;
wire \op2[8] ;
wire \op2[7] ;
wire \op2[6] ;
wire \op2[5] ;
wire \op2[4] ;
wire \op2[3] ;
wire \op2[2] ;
wire \op2[1] ;
wire \op1[31] ;
wire \op1[30] ;
wire \op1[29] ;
wire \op1[28] ;
wire \op1[27] ;
wire \op1[26] ;
wire \op1[25] ;
wire \op1[24] ;
wire \op1[23] ;
wire \op1[22] ;
wire \op1[21] ;
wire \op1[20] ;
wire \op1[19] ;
wire \op1[18] ;
wire \op1[17] ;
wire \op1[16] ;
wire \op1[15] ;
wire \op1[14] ;
wire \op1[13] ;
wire \op1[12] ;
wire \op1[11] ;
wire \op1[10] ;
wire \op1[9] ;
wire \op1[8] ;
wire \op1[7] ;
wire \op1[6] ;
wire \op1[5] ;
wire \op1[4] ;
wire \op1[3] ;
wire \op1[2] ;
wire \op1[1] ;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_1_7;
wire n_0_1_8;
wire n_0_1_9;
wire n_0_1_10;
wire n_0_1_12;
wire hfn_ipo_n7;
wire n_0_1_14;
wire n_0_1_15;
wire n_0_1_16;
wire n_0_1_17;
wire n_0_1_18;
wire n_0_1_19;
wire n_0_1_20;
wire n_0_1_21;
wire n_0_1_22;
wire n_0_1_23;
wire n_0_1_24;
wire n_0_1_25;
wire n_0_1_26;
wire n_0_1_27;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_1_30;
wire hfn_ipo_n8;
wire n_0_1_1;
wire n_0_1_2;
wire n_0_1_3;
wire n_0_1_4;
wire n_0_1_11;
wire uc_0;
wire uc_1;
wire uc_2;
wire n_0;
wire uc_3;
wire uc_4;
wire uc_5;
wire n_1;
wire uc_6;
wire uc_7;
wire uc_8;
wire n_2;
wire uc_9;
wire uc_10;
wire uc_11;
wire n_3;
wire uc_12;
wire uc_13;
wire uc_14;
wire n_4;
wire uc_15;
wire uc_16;
wire uc_17;
wire n_5;
wire uc_18;
wire uc_19;
wire uc_20;
wire n_6;
wire uc_21;
wire uc_22;
wire uc_23;
wire n_7;
wire uc_24;
wire uc_25;
wire uc_26;
wire n_8;
wire uc_27;
wire uc_28;
wire uc_29;
wire n_9;
wire uc_30;
wire uc_31;
wire uc_32;
wire n_10;
wire uc_33;
wire uc_34;
wire uc_35;
wire n_11;
wire uc_36;
wire uc_37;
wire uc_38;
wire n_12;
wire uc_39;
wire uc_40;
wire uc_41;
wire n_13;
wire uc_42;
wire uc_43;
wire uc_44;
wire n_14;
wire uc_45;
wire uc_46;
wire uc_47;
wire n_15;
wire uc_48;
wire uc_49;
wire uc_50;
wire n_16;
wire uc_51;
wire uc_52;
wire uc_53;
wire n_17;
wire uc_54;
wire uc_55;
wire uc_56;
wire n_18;
wire uc_57;
wire uc_58;
wire uc_59;
wire n_19;
wire uc_60;
wire uc_61;
wire uc_62;
wire n_20;
wire uc_63;
wire uc_64;
wire uc_65;
wire n_21;
wire uc_66;
wire uc_67;
wire uc_68;
wire n_22;
wire uc_69;
wire uc_70;
wire uc_71;
wire n_23;
wire uc_72;
wire uc_73;
wire uc_74;
wire n_24;
wire uc_75;
wire uc_76;
wire uc_77;
wire n_25;
wire uc_78;
wire uc_79;
wire uc_80;
wire n_26;
wire uc_81;
wire uc_82;
wire uc_83;
wire n_27;
wire uc_84;
wire uc_85;
wire uc_86;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;


XNOR2_X1 i_0_1_155 (.ZN (n_0_1_11), .A (b[31]), .B (a[31]));
NAND2_X1 i_0_1_154 (.ZN (n_0_1_4), .A1 (n_55), .A2 (hfn_ipo_n8));
NAND2_X1 i_0_1_153 (.ZN (n_0_1_3), .A1 (n_0_1_12), .A2 (a[22]));
NAND2_X1 i_0_1_152 (.ZN (n_0_1_2), .A1 (n_0_21), .A2 (a[31]));
NAND2_X2 i_0_1_151 (.ZN (\op1[22] ), .A1 (n_0_1_2), .A2 (n_0_1_3));
NAND2_X1 i_0_1_150 (.ZN (n_0_1_1), .A1 (a[31]), .A2 (n_0_26));
CLKBUF_X1 hfn_ipo_c8 (.Z (hfn_ipo_n8), .A (n_0_1_11));
NAND2_X1 i_0_1_148 (.ZN (n_0_1_30), .A1 (n_0_1_12), .A2 (a[27]));
NAND2_X1 i_0_1_147 (.ZN (\op1[27] ), .A1 (n_0_1_30), .A2 (n_0_1_1));
NAND2_X1 i_0_1_146 (.ZN (n_0_1_29), .A1 (a[31]), .A2 (n_0_25));
NAND2_X1 i_0_1_145 (.ZN (n_0_1_28), .A1 (n_0_1_12), .A2 (a[26]));
NAND2_X2 i_0_1_144 (.ZN (\op1[26] ), .A1 (n_0_1_28), .A2 (n_0_1_29));
NAND2_X1 i_0_1_143 (.ZN (n_0_1_27), .A1 (a[31]), .A2 (n_0_24));
NAND2_X1 i_0_1_142 (.ZN (n_0_1_26), .A1 (n_0_1_12), .A2 (a[25]));
NAND2_X2 i_0_1_141 (.ZN (\op1[25] ), .A1 (n_0_1_26), .A2 (n_0_1_27));
NAND2_X1 i_0_1_140 (.ZN (n_0_1_25), .A1 (a[31]), .A2 (n_0_23));
NAND2_X1 i_0_1_139 (.ZN (n_0_1_24), .A1 (a[24]), .A2 (n_0_1_12));
NAND2_X2 i_0_1_138 (.ZN (\op1[24] ), .A1 (n_0_1_25), .A2 (n_0_1_24));
NAND2_X1 i_0_1_137 (.ZN (n_0_1_23), .A1 (a[31]), .A2 (n_0_22));
NAND2_X1 i_0_1_136 (.ZN (n_0_1_22), .A1 (n_0_1_12), .A2 (a[23]));
NAND2_X1 i_0_1_135 (.ZN (\op1[23] ), .A1 (n_0_1_22), .A2 (n_0_1_23));
NAND2_X1 i_0_1_134 (.ZN (n_0_1_21), .A1 (a[31]), .A2 (n_0_20));
NAND2_X1 i_0_1_133 (.ZN (n_0_1_20), .A1 (n_0_1_12), .A2 (a[21]));
NAND2_X1 i_0_1_132 (.ZN (\op1[21] ), .A1 (n_0_1_20), .A2 (n_0_1_21));
NAND2_X1 i_0_1_131 (.ZN (n_0_1_19), .A1 (a[31]), .A2 (n_0_19));
NAND2_X1 i_0_1_130 (.ZN (n_0_1_18), .A1 (a[20]), .A2 (n_0_1_12));
NAND2_X2 i_0_1_129 (.ZN (\op1[20] ), .A1 (n_0_1_19), .A2 (n_0_1_18));
NAND2_X1 i_0_1_128 (.ZN (n_0_1_17), .A1 (a[31]), .A2 (n_0_18));
NAND2_X1 i_0_1_123 (.ZN (n_0_1_16), .A1 (n_0_1_12), .A2 (a[19]));
NAND2_X1 i_0_1_122 (.ZN (\op1[19] ), .A1 (n_0_1_16), .A2 (n_0_1_17));
NAND2_X1 i_0_1_121 (.ZN (n_0_1_15), .A1 (a[31]), .A2 (n_0_17));
NAND2_X1 i_0_1_120 (.ZN (n_0_1_14), .A1 (n_0_1_12), .A2 (a[18]));
NAND2_X1 i_0_1_119 (.ZN (\op1[18] ), .A1 (n_0_1_14), .A2 (n_0_1_15));
CLKBUF_X3 hfn_ipo_c7 (.Z (hfn_ipo_n7), .A (n_0_1_11));
INV_X1 i_0_1_57 (.ZN (n_0_1_12), .A (a[31]));
INV_X1 i_0_1_56 (.ZN (n_0_1_10), .A (hfn_ipo_n8));
NAND2_X1 i_0_1_55 (.ZN (n_0_1_9), .A1 (n_0_124), .A2 (n_0_1_10));
NAND2_X1 i_0_1_54 (.ZN (n_0_1_8), .A1 (n_28), .A2 (hfn_ipo_n8));
NAND2_X1 i_0_1_53 (.ZN (out[63]), .A1 (n_0_1_9), .A2 (n_0_1_8));
INV_X1 i_0_1_52 (.ZN (n_0_1_7), .A (n_0_123));
NAND2_X1 i_0_1_51 (.ZN (n_0_1_6), .A1 (n_60), .A2 (hfn_ipo_n8));
OAI21_X1 i_0_1_50 (.ZN (out[62]), .A (n_0_1_6), .B1 (n_0_1_7), .B2 (hfn_ipo_n8));
MUX2_X1 i_0_1_127 (.Z (out[61]), .A (n_0_122), .B (n_59), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_126 (.Z (out[60]), .A (n_0_121), .B (n_58), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_125 (.Z (out[59]), .A (n_0_120), .B (n_57), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_124 (.Z (out[58]), .A (n_0_119), .B (n_56), .S (hfn_ipo_n8));
INV_X1 i_0_1_49 (.ZN (n_0_1_5), .A (n_0_118));
OAI21_X1 i_0_1_0 (.ZN (out[57]), .A (n_0_1_4), .B1 (n_0_1_5), .B2 (hfn_ipo_n8));
MUX2_X1 i_0_1_118 (.Z (out[56]), .A (n_0_117), .B (n_54), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_117 (.Z (out[55]), .A (n_0_116), .B (n_53), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_116 (.Z (out[54]), .A (n_0_115), .B (n_52), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_115 (.Z (out[53]), .A (n_0_114), .B (n_51), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_114 (.Z (out[52]), .A (n_0_113), .B (n_50), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_113 (.Z (out[51]), .A (n_0_112), .B (n_49), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_112 (.Z (out[50]), .A (n_0_111), .B (n_48), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_111 (.Z (out[49]), .A (n_0_110), .B (n_47), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_110 (.Z (out[48]), .A (n_0_109), .B (n_46), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_109 (.Z (out[47]), .A (n_0_108), .B (n_45), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_108 (.Z (out[46]), .A (n_0_107), .B (n_44), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_107 (.Z (out[45]), .A (n_0_106), .B (n_43), .S (hfn_ipo_n8));
MUX2_X1 i_0_1_106 (.Z (out[44]), .A (n_0_105), .B (n_42), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_105 (.Z (out[43]), .A (n_0_104), .B (n_41), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_104 (.Z (out[42]), .A (n_0_103), .B (n_40), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_103 (.Z (out[41]), .A (n_0_102), .B (n_39), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_102 (.Z (out[40]), .A (n_0_101), .B (n_38), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_101 (.Z (out[39]), .A (n_0_100), .B (n_37), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_100 (.Z (out[38]), .A (n_0_99), .B (n_36), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_99 (.Z (out[37]), .A (n_0_98), .B (n_35), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_98 (.Z (out[36]), .A (n_0_97), .B (n_34), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_97 (.Z (out[35]), .A (n_0_96), .B (n_33), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_96 (.Z (out[34]), .A (n_0_95), .B (n_32), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_95 (.Z (out[33]), .A (n_0_94), .B (n_31), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_94 (.Z (out[32]), .A (n_0_93), .B (n_30), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_93 (.Z (out[31]), .A (n_0_92), .B (n_29), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_92 (.Z (out[30]), .A (n_0_91), .B (\s1[29][0] ), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_91 (.Z (out[29]), .A (n_0_90), .B (n_27), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_90 (.Z (out[28]), .A (n_0_89), .B (n_26), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_89 (.Z (out[27]), .A (n_0_88), .B (n_25), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_88 (.Z (out[26]), .A (n_0_87), .B (n_24), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_87 (.Z (out[25]), .A (n_0_86), .B (n_23), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_86 (.Z (out[24]), .A (n_0_85), .B (n_22), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_85 (.Z (out[23]), .A (n_0_84), .B (n_21), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_84 (.Z (out[22]), .A (n_0_83), .B (n_20), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_83 (.Z (out[21]), .A (n_0_82), .B (n_19), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_82 (.Z (out[20]), .A (n_0_81), .B (n_18), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_81 (.Z (out[19]), .A (n_0_80), .B (n_17), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_80 (.Z (out[18]), .A (n_0_79), .B (n_16), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_79 (.Z (out[17]), .A (n_0_78), .B (n_15), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_78 (.Z (out[16]), .A (n_0_77), .B (n_14), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_77 (.Z (out[15]), .A (n_0_76), .B (n_13), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_76 (.Z (out[14]), .A (n_0_75), .B (n_12), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_75 (.Z (out[13]), .A (n_0_74), .B (n_11), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_74 (.Z (out[12]), .A (n_0_73), .B (n_10), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_73 (.Z (out[11]), .A (n_0_72), .B (n_9), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_72 (.Z (out[10]), .A (n_0_71), .B (n_8), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_71 (.Z (out[9]), .A (n_0_70), .B (n_7), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_70 (.Z (out[8]), .A (n_0_69), .B (n_6), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_69 (.Z (out[7]), .A (n_0_68), .B (n_5), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_68 (.Z (out[6]), .A (n_0_67), .B (n_4), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_67 (.Z (out[5]), .A (n_0_66), .B (n_3), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_66 (.Z (out[4]), .A (n_0_65), .B (n_2), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_65 (.Z (out[3]), .A (n_0_64), .B (n_1), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_64 (.Z (out[2]), .A (n_0_63), .B (n_0), .S (hfn_ipo_n7));
MUX2_X1 i_0_1_63 (.Z (out[1]), .A (n_0_62), .B (\s1[0][0] ), .S (hfn_ipo_n7));
AND2_X1 i_0_1_62 (.ZN (\op1[31] ), .A1 (n_0_30), .A2 (a[31]));
MUX2_X1 i_0_1_61 (.Z (\op1[30] ), .A (a[30]), .B (n_0_29), .S (a[31]));
MUX2_X1 i_0_1_60 (.Z (\op1[29] ), .A (a[29]), .B (n_0_28), .S (a[31]));
MUX2_X1 i_0_1_59 (.Z (\op1[28] ), .A (a[28]), .B (n_0_27), .S (a[31]));
MUX2_X1 i_0_1_48 (.Z (\op1[17] ), .A (a[17]), .B (n_0_16), .S (a[31]));
MUX2_X1 i_0_1_47 (.Z (\op1[16] ), .A (a[16]), .B (n_0_15), .S (a[31]));
MUX2_X1 i_0_1_46 (.Z (\op1[15] ), .A (a[15]), .B (n_0_14), .S (a[31]));
MUX2_X1 i_0_1_45 (.Z (\op1[14] ), .A (a[14]), .B (n_0_13), .S (a[31]));
MUX2_X1 i_0_1_44 (.Z (\op1[13] ), .A (a[13]), .B (n_0_12), .S (a[31]));
MUX2_X1 i_0_1_43 (.Z (\op1[12] ), .A (a[12]), .B (n_0_11), .S (a[31]));
MUX2_X1 i_0_1_42 (.Z (\op1[11] ), .A (a[11]), .B (n_0_10), .S (a[31]));
MUX2_X1 i_0_1_41 (.Z (\op1[10] ), .A (a[10]), .B (n_0_9), .S (a[31]));
MUX2_X1 i_0_1_40 (.Z (\op1[9] ), .A (a[9]), .B (n_0_8), .S (a[31]));
MUX2_X1 i_0_1_39 (.Z (\op1[8] ), .A (a[8]), .B (n_0_7), .S (a[31]));
MUX2_X1 i_0_1_38 (.Z (\op1[7] ), .A (a[7]), .B (n_0_6), .S (a[31]));
MUX2_X1 i_0_1_37 (.Z (\op1[6] ), .A (a[6]), .B (n_0_5), .S (a[31]));
MUX2_X1 i_0_1_36 (.Z (\op1[5] ), .A (a[5]), .B (n_0_4), .S (a[31]));
MUX2_X1 i_0_1_35 (.Z (\op1[4] ), .A (a[4]), .B (n_0_3), .S (a[31]));
MUX2_X1 i_0_1_34 (.Z (\op1[3] ), .A (a[3]), .B (n_0_2), .S (a[31]));
MUX2_X1 i_0_1_33 (.Z (\op1[2] ), .A (a[2]), .B (n_0_1), .S (a[31]));
MUX2_X1 i_0_1_32 (.Z (\op1[1] ), .A (a[1]), .B (n_0_0), .S (a[31]));
AND2_X1 i_0_1_31 (.ZN (\op2[31] ), .A1 (n_0_61), .A2 (b[31]));
MUX2_X1 i_0_1_30 (.Z (\op2[30] ), .A (b[30]), .B (n_0_60), .S (b[31]));
MUX2_X1 i_0_1_29 (.Z (\op2[29] ), .A (b[29]), .B (n_0_59), .S (b[31]));
MUX2_X1 i_0_1_28 (.Z (\op2[28] ), .A (b[28]), .B (n_0_58), .S (b[31]));
MUX2_X1 i_0_1_27 (.Z (\op2[27] ), .A (b[27]), .B (n_0_57), .S (b[31]));
MUX2_X1 i_0_1_26 (.Z (\op2[26] ), .A (b[26]), .B (n_0_56), .S (b[31]));
MUX2_X1 i_0_1_25 (.Z (\op2[25] ), .A (b[25]), .B (n_0_55), .S (b[31]));
MUX2_X1 i_0_1_24 (.Z (\op2[24] ), .A (b[24]), .B (n_0_54), .S (b[31]));
MUX2_X1 i_0_1_23 (.Z (\op2[23] ), .A (b[23]), .B (n_0_53), .S (b[31]));
MUX2_X1 i_0_1_22 (.Z (\op2[22] ), .A (b[22]), .B (n_0_52), .S (b[31]));
MUX2_X1 i_0_1_21 (.Z (\op2[21] ), .A (b[21]), .B (n_0_51), .S (b[31]));
MUX2_X1 i_0_1_20 (.Z (\op2[20] ), .A (b[20]), .B (n_0_50), .S (b[31]));
MUX2_X1 i_0_1_19 (.Z (\op2[19] ), .A (b[19]), .B (n_0_49), .S (b[31]));
MUX2_X1 i_0_1_18 (.Z (\op2[18] ), .A (b[18]), .B (n_0_48), .S (b[31]));
MUX2_X1 i_0_1_17 (.Z (\op2[17] ), .A (b[17]), .B (n_0_47), .S (b[31]));
MUX2_X1 i_0_1_16 (.Z (\op2[16] ), .A (b[16]), .B (n_0_46), .S (b[31]));
MUX2_X1 i_0_1_15 (.Z (\op2[15] ), .A (b[15]), .B (n_0_45), .S (b[31]));
MUX2_X1 i_0_1_14 (.Z (\op2[14] ), .A (b[14]), .B (n_0_44), .S (b[31]));
MUX2_X1 i_0_1_13 (.Z (\op2[13] ), .A (b[13]), .B (n_0_43), .S (b[31]));
MUX2_X1 i_0_1_12 (.Z (\op2[12] ), .A (b[12]), .B (n_0_42), .S (b[31]));
MUX2_X1 i_0_1_11 (.Z (\op2[11] ), .A (b[11]), .B (n_0_41), .S (b[31]));
MUX2_X1 i_0_1_10 (.Z (\op2[10] ), .A (b[10]), .B (n_0_40), .S (b[31]));
MUX2_X1 i_0_1_9 (.Z (\op2[9] ), .A (b[9]), .B (n_0_39), .S (b[31]));
MUX2_X1 i_0_1_8 (.Z (\op2[8] ), .A (b[8]), .B (n_0_38), .S (b[31]));
MUX2_X1 i_0_1_7 (.Z (\op2[7] ), .A (b[7]), .B (n_0_37), .S (b[31]));
MUX2_X1 i_0_1_6 (.Z (\op2[6] ), .A (b[6]), .B (n_0_36), .S (b[31]));
MUX2_X1 i_0_1_5 (.Z (\op2[5] ), .A (b[5]), .B (n_0_35), .S (b[31]));
MUX2_X1 i_0_1_4 (.Z (\op2[4] ), .A (b[4]), .B (n_0_34), .S (b[31]));
MUX2_X1 i_0_1_3 (.Z (\op2[3] ), .A (b[3]), .B (n_0_33), .S (b[31]));
MUX2_X1 i_0_1_2 (.Z (\op2[2] ), .A (b[2]), .B (n_0_32), .S (b[31]));
MUX2_X1 i_0_1_1 (.Z (\op2[1] ), .A (b[1]), .B (n_0_31), .S (b[31]));
datapath__0_38 i_0_36 (.p_0 ({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, 
    n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
    n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
    n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
    n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
    n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
    n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, uc_93})
    , .sum1 ({n_28, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
    n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, \s1[29][0] , n_27, n_26, n_25, 
    n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, \s1[0][0] , out[0]}));
datapath__0_3 i_0_0 (.p_0 ({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
    n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
    n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
    n_0_2, n_0_1, n_0_0, uc_92}), .a ({a[31], a[30], a[29], a[28], a[27], a[26], 
    a[25], a[24], a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16], a[15], 
    a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], 
    a[2], a[1], a[0]}));
datapath__0_4 i_0_2 (.p_0 ({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
    n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
    n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
    n_0_34, n_0_33, n_0_32, n_0_31, uc_91}), .b ({b[31], b[30], b[29], b[28], b[27], 
    b[26], b[25], b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], 
    b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], 
    b[3], b[2], b[1], b[0]}));
PartialAdder p1 (.c1 ({\c1[0][31] , \c1[0][30] , \c1[0][29] , \c1[0][28] , \c1[0][27] , 
    \c1[0][26] , \c1[0][25] , \c1[0][24] , \c1[0][23] , \c1[0][22] , \c1[0][21] , 
    \c1[0][20] , \c1[0][19] , \c1[0][18] , \c1[0][17] , \c1[0][16] , \c1[0][15] , 
    \c1[0][14] , \c1[0][13] , \c1[0][12] , \c1[0][11] , \c1[0][10] , \c1[0][9] , 
    \c1[0][8] , \c1[0][7] , \c1[0][6] , \c1[0][5] , \c1[0][4] , \c1[0][3] , \c1[0][2] , 
    \c1[0][1] , \c1[0][0] }), .s1 ({uc_90, \s1[0][31] , \s1[0][30] , \s1[0][29] , 
    \s1[0][28] , \s1[0][27] , \s1[0][26] , \s1[0][25] , \s1[0][24] , \s1[0][23] , 
    \s1[0][22] , \s1[0][21] , \s1[0][20] , \s1[0][19] , \s1[0][18] , \s1[0][17] , 
    \s1[0][16] , \s1[0][15] , \s1[0][14] , \s1[0][13] , \s1[0][12] , \s1[0][11] , 
    \s1[0][10] , \s1[0][9] , \s1[0][8] , \s1[0][7] , \s1[0][6] , \s1[0][5] , \s1[0][4] , 
    \s1[0][3] , \s1[0][2] , \s1[0][1] , \s1[0][0] }), .a ({uc_87, \partial_reg[0][31] , 
    \partial_reg[0][30] , \partial_reg[0][29] , \partial_reg[0][28] , \partial_reg[0][27] , 
    \partial_reg[0][26] , \partial_reg[0][25] , \partial_reg[0][24] , \partial_reg[0][23] , 
    \partial_reg[0][22] , \partial_reg[0][21] , \partial_reg[0][20] , \partial_reg[0][19] , 
    \partial_reg[0][18] , \partial_reg[0][17] , \partial_reg[0][16] , \partial_reg[0][15] , 
    \partial_reg[0][14] , \partial_reg[0][13] , \partial_reg[0][12] , \partial_reg[0][11] , 
    \partial_reg[0][10] , \partial_reg[0][9] , \partial_reg[0][8] , \partial_reg[0][7] , 
    \partial_reg[0][6] , \partial_reg[0][5] , \partial_reg[0][4] , \partial_reg[0][3] , 
    \partial_reg[0][2] , \partial_reg[0][1] , uc_88}), .b ({\partial_reg[1][31] , 
    \partial_reg[1][30] , \partial_reg[1][29] , \partial_reg[1][28] , \partial_reg[1][27] , 
    \partial_reg[1][26] , \partial_reg[1][25] , \partial_reg[1][24] , \partial_reg[1][23] , 
    \partial_reg[1][22] , \partial_reg[1][21] , \partial_reg[1][20] , \partial_reg[1][19] , 
    \partial_reg[1][18] , \partial_reg[1][17] , \partial_reg[1][16] , \partial_reg[1][15] , 
    \partial_reg[1][14] , \partial_reg[1][13] , \partial_reg[1][12] , \partial_reg[1][11] , 
    \partial_reg[1][10] , \partial_reg[1][9] , \partial_reg[1][8] , \partial_reg[1][7] , 
    \partial_reg[1][6] , \partial_reg[1][5] , \partial_reg[1][4] , \partial_reg[1][3] , 
    \partial_reg[1][2] , \partial_reg[1][1] , \partial_reg[1][0] }), .c ({uc_89, 
    \partial_reg[2][30] , \partial_reg[2][29] , \partial_reg[2][28] , \partial_reg[2][27] , 
    \partial_reg[2][26] , \partial_reg[2][25] , \partial_reg[2][24] , \partial_reg[2][23] , 
    \partial_reg[2][22] , \partial_reg[2][21] , \partial_reg[2][20] , \partial_reg[2][19] , 
    \partial_reg[2][18] , \partial_reg[2][17] , \partial_reg[2][16] , \partial_reg[2][15] , 
    \partial_reg[2][14] , \partial_reg[2][13] , \partial_reg[2][12] , \partial_reg[2][11] , 
    \partial_reg[2][10] , \partial_reg[2][9] , \partial_reg[2][8] , \partial_reg[2][7] , 
    \partial_reg[2][6] , \partial_reg[2][5] , \partial_reg[2][4] , \partial_reg[2][3] , 
    \partial_reg[2][2] , \partial_reg[2][1] , \partial_reg[2][0] }));
AND2_X1 i_4_0_1089 (.ZN (\partial_reg[2][30] ), .A1 (\op1[30] ), .A2 (\op2[2] ));
AND2_X1 i_4_0_1088 (.ZN (\partial_reg[2][29] ), .A1 (\op1[29] ), .A2 (\op2[2] ));
AND2_X1 i_4_0_129 (.ZN (\partial_reg[0][31] ), .A1 (\op1[31] ), .A2 (b[0]));
NAND2_X1 i_4_0_128 (.ZN (n_4_0_65), .A1 (\op1[31] ), .A2 (\op2[1] ));
INV_X1 i_4_0_98 (.ZN (\partial_reg[1][31] ), .A (n_4_0_65));
NAND2_X1 i_4_0_97 (.ZN (n_4_0_64), .A1 (\op1[30] ), .A2 (\op2[1] ));
INV_X1 i_4_0_96 (.ZN (\partial_reg[1][30] ), .A (n_4_0_64));
INV_X2 i_4_0_65 (.ZN (n_4_0_0), .A (b[0]));
INV_X2 i_4_0_64 (.ZN (n_4_0_30), .A (\op1[29] ));
INV_X2 i_4_0_63 (.ZN (n_4_0_31), .A (\op1[30] ));
INV_X2 i_4_0_61 (.ZN (n_4_0_32), .A (\op1[31] ));
INV_X2 i_4_0_59 (.ZN (n_4_0_33), .A (\op2[1] ));
INV_X4 i_4_0_0 (.ZN (n_4_0_34), .A (\op2[2] ));
NOR2_X1 i_4_0_1087 (.ZN (\partial_reg[31][31] ), .A1 (n_4_0_32), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1086 (.ZN (\partial_reg[31][30] ), .A1 (n_4_0_31), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1085 (.ZN (\partial_reg[31][29] ), .A1 (n_4_0_30), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1084 (.ZN (\partial_reg[31][28] ), .A1 (n_4_0_29), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1083 (.ZN (\partial_reg[31][27] ), .A1 (n_4_0_28), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1082 (.ZN (\partial_reg[31][26] ), .A1 (n_4_0_27), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1081 (.ZN (\partial_reg[31][25] ), .A1 (n_4_0_26), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1080 (.ZN (\partial_reg[31][24] ), .A1 (n_4_0_25), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1079 (.ZN (\partial_reg[31][23] ), .A1 (n_4_0_24), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1078 (.ZN (\partial_reg[31][22] ), .A1 (n_4_0_23), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1077 (.ZN (\partial_reg[31][21] ), .A1 (n_4_0_22), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1076 (.ZN (\partial_reg[31][20] ), .A1 (n_4_0_21), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1075 (.ZN (\partial_reg[31][19] ), .A1 (n_4_0_20), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1074 (.ZN (\partial_reg[31][18] ), .A1 (n_4_0_19), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1073 (.ZN (\partial_reg[31][17] ), .A1 (n_4_0_18), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1072 (.ZN (\partial_reg[31][16] ), .A1 (n_4_0_17), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1071 (.ZN (\partial_reg[31][15] ), .A1 (n_4_0_16), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1070 (.ZN (\partial_reg[31][14] ), .A1 (n_4_0_15), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1069 (.ZN (\partial_reg[31][13] ), .A1 (n_4_0_14), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1068 (.ZN (\partial_reg[31][12] ), .A1 (n_4_0_13), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1067 (.ZN (\partial_reg[31][11] ), .A1 (n_4_0_12), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1066 (.ZN (\partial_reg[31][10] ), .A1 (n_4_0_11), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1065 (.ZN (\partial_reg[31][9] ), .A1 (n_4_0_10), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1064 (.ZN (\partial_reg[31][8] ), .A1 (n_4_0_9), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1063 (.ZN (\partial_reg[31][7] ), .A1 (n_4_0_8), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1062 (.ZN (\partial_reg[31][6] ), .A1 (n_4_0_7), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1061 (.ZN (\partial_reg[31][5] ), .A1 (n_4_0_6), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1060 (.ZN (\partial_reg[31][4] ), .A1 (n_4_0_5), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1059 (.ZN (\partial_reg[31][3] ), .A1 (n_4_0_4), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1058 (.ZN (\partial_reg[31][2] ), .A1 (n_4_0_3), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1057 (.ZN (\partial_reg[31][1] ), .A1 (n_4_0_2), .A2 (n_4_0_63));
NOR2_X1 i_4_0_1056 (.ZN (\partial_reg[31][0] ), .A1 (n_4_0_1), .A2 (n_4_0_63));
INV_X2 i_4_0_1055 (.ZN (n_4_0_63), .A (\op2[31] ));
NOR2_X1 i_4_0_1054 (.ZN (\partial_reg[30][31] ), .A1 (n_4_0_62), .A2 (n_4_0_32));
NOR2_X1 i_4_0_1053 (.ZN (\partial_reg[30][30] ), .A1 (n_4_0_62), .A2 (n_4_0_31));
NOR2_X1 i_4_0_1052 (.ZN (\partial_reg[30][29] ), .A1 (n_4_0_62), .A2 (n_4_0_30));
NOR2_X1 i_4_0_1051 (.ZN (\partial_reg[30][28] ), .A1 (n_4_0_62), .A2 (n_4_0_29));
NOR2_X1 i_4_0_1050 (.ZN (\partial_reg[30][27] ), .A1 (n_4_0_62), .A2 (n_4_0_28));
NOR2_X1 i_4_0_1049 (.ZN (\partial_reg[30][26] ), .A1 (n_4_0_62), .A2 (n_4_0_27));
NOR2_X1 i_4_0_1048 (.ZN (\partial_reg[30][25] ), .A1 (n_4_0_62), .A2 (n_4_0_26));
NOR2_X1 i_4_0_1047 (.ZN (\partial_reg[30][24] ), .A1 (n_4_0_62), .A2 (n_4_0_25));
NOR2_X1 i_4_0_1046 (.ZN (\partial_reg[30][23] ), .A1 (n_4_0_62), .A2 (n_4_0_24));
NOR2_X1 i_4_0_1045 (.ZN (\partial_reg[30][22] ), .A1 (n_4_0_62), .A2 (n_4_0_23));
NOR2_X1 i_4_0_1044 (.ZN (\partial_reg[30][21] ), .A1 (n_4_0_62), .A2 (n_4_0_22));
NOR2_X1 i_4_0_1043 (.ZN (\partial_reg[30][20] ), .A1 (n_4_0_62), .A2 (n_4_0_21));
NOR2_X1 i_4_0_1042 (.ZN (\partial_reg[30][19] ), .A1 (n_4_0_62), .A2 (n_4_0_20));
NOR2_X1 i_4_0_1041 (.ZN (\partial_reg[30][18] ), .A1 (n_4_0_62), .A2 (n_4_0_19));
NOR2_X1 i_4_0_1040 (.ZN (\partial_reg[30][17] ), .A1 (n_4_0_62), .A2 (n_4_0_18));
NOR2_X1 i_4_0_1039 (.ZN (\partial_reg[30][16] ), .A1 (n_4_0_62), .A2 (n_4_0_17));
NOR2_X1 i_4_0_1038 (.ZN (\partial_reg[30][15] ), .A1 (n_4_0_62), .A2 (n_4_0_16));
NOR2_X1 i_4_0_1037 (.ZN (\partial_reg[30][14] ), .A1 (n_4_0_62), .A2 (n_4_0_15));
NOR2_X1 i_4_0_1036 (.ZN (\partial_reg[30][13] ), .A1 (n_4_0_62), .A2 (n_4_0_14));
NOR2_X1 i_4_0_1035 (.ZN (\partial_reg[30][12] ), .A1 (n_4_0_62), .A2 (n_4_0_13));
NOR2_X1 i_4_0_1034 (.ZN (\partial_reg[30][11] ), .A1 (n_4_0_62), .A2 (n_4_0_12));
NOR2_X1 i_4_0_1033 (.ZN (\partial_reg[30][10] ), .A1 (n_4_0_62), .A2 (n_4_0_11));
NOR2_X1 i_4_0_1032 (.ZN (\partial_reg[30][9] ), .A1 (n_4_0_62), .A2 (n_4_0_10));
NOR2_X1 i_4_0_1031 (.ZN (\partial_reg[30][8] ), .A1 (n_4_0_62), .A2 (n_4_0_9));
NOR2_X1 i_4_0_1030 (.ZN (\partial_reg[30][7] ), .A1 (n_4_0_62), .A2 (n_4_0_8));
NOR2_X1 i_4_0_1029 (.ZN (\partial_reg[30][6] ), .A1 (n_4_0_62), .A2 (n_4_0_7));
NOR2_X1 i_4_0_1028 (.ZN (\partial_reg[30][5] ), .A1 (n_4_0_62), .A2 (n_4_0_6));
NOR2_X1 i_4_0_1027 (.ZN (\partial_reg[30][4] ), .A1 (n_4_0_62), .A2 (n_4_0_5));
NOR2_X1 i_4_0_1026 (.ZN (\partial_reg[30][3] ), .A1 (n_4_0_62), .A2 (n_4_0_4));
NOR2_X1 i_4_0_1025 (.ZN (\partial_reg[30][2] ), .A1 (n_4_0_62), .A2 (n_4_0_3));
NOR2_X1 i_4_0_1024 (.ZN (\partial_reg[30][1] ), .A1 (n_4_0_62), .A2 (n_4_0_2));
NOR2_X2 i_4_0_1023 (.ZN (\partial_reg[30][0] ), .A1 (n_4_0_62), .A2 (n_4_0_1));
INV_X2 i_4_0_1022 (.ZN (n_4_0_62), .A (\op2[30] ));
NOR2_X1 i_4_0_1021 (.ZN (\partial_reg[29][31] ), .A1 (n_4_0_61), .A2 (n_4_0_32));
NOR2_X1 i_4_0_1020 (.ZN (\partial_reg[29][30] ), .A1 (n_4_0_61), .A2 (n_4_0_31));
NOR2_X1 i_4_0_1019 (.ZN (\partial_reg[29][29] ), .A1 (n_4_0_61), .A2 (n_4_0_30));
NOR2_X1 i_4_0_1018 (.ZN (\partial_reg[29][28] ), .A1 (n_4_0_61), .A2 (n_4_0_29));
NOR2_X1 i_4_0_1017 (.ZN (\partial_reg[29][27] ), .A1 (n_4_0_61), .A2 (n_4_0_28));
NOR2_X1 i_4_0_1016 (.ZN (\partial_reg[29][26] ), .A1 (n_4_0_61), .A2 (n_4_0_27));
NOR2_X1 i_4_0_1015 (.ZN (\partial_reg[29][25] ), .A1 (n_4_0_61), .A2 (n_4_0_26));
NOR2_X1 i_4_0_1014 (.ZN (\partial_reg[29][24] ), .A1 (n_4_0_61), .A2 (n_4_0_25));
NOR2_X1 i_4_0_1013 (.ZN (\partial_reg[29][23] ), .A1 (n_4_0_61), .A2 (n_4_0_24));
NOR2_X1 i_4_0_1012 (.ZN (\partial_reg[29][22] ), .A1 (n_4_0_61), .A2 (n_4_0_23));
NOR2_X1 i_4_0_1011 (.ZN (\partial_reg[29][21] ), .A1 (n_4_0_61), .A2 (n_4_0_22));
NOR2_X1 i_4_0_1010 (.ZN (\partial_reg[29][20] ), .A1 (n_4_0_61), .A2 (n_4_0_21));
NOR2_X1 i_4_0_1009 (.ZN (\partial_reg[29][19] ), .A1 (n_4_0_61), .A2 (n_4_0_20));
NOR2_X1 i_4_0_1008 (.ZN (\partial_reg[29][18] ), .A1 (n_4_0_61), .A2 (n_4_0_19));
NOR2_X1 i_4_0_1007 (.ZN (\partial_reg[29][17] ), .A1 (n_4_0_61), .A2 (n_4_0_18));
NOR2_X1 i_4_0_1006 (.ZN (\partial_reg[29][16] ), .A1 (n_4_0_61), .A2 (n_4_0_17));
NOR2_X1 i_4_0_1005 (.ZN (\partial_reg[29][15] ), .A1 (n_4_0_61), .A2 (n_4_0_16));
NOR2_X1 i_4_0_1004 (.ZN (\partial_reg[29][14] ), .A1 (n_4_0_61), .A2 (n_4_0_15));
NOR2_X1 i_4_0_1003 (.ZN (\partial_reg[29][13] ), .A1 (n_4_0_61), .A2 (n_4_0_14));
NOR2_X1 i_4_0_1002 (.ZN (\partial_reg[29][12] ), .A1 (n_4_0_61), .A2 (n_4_0_13));
NOR2_X1 i_4_0_1001 (.ZN (\partial_reg[29][11] ), .A1 (n_4_0_61), .A2 (n_4_0_12));
NOR2_X1 i_4_0_1000 (.ZN (\partial_reg[29][10] ), .A1 (n_4_0_61), .A2 (n_4_0_11));
NOR2_X1 i_4_0_999 (.ZN (\partial_reg[29][9] ), .A1 (n_4_0_61), .A2 (n_4_0_10));
NOR2_X1 i_4_0_998 (.ZN (\partial_reg[29][8] ), .A1 (n_4_0_61), .A2 (n_4_0_9));
NOR2_X1 i_4_0_997 (.ZN (\partial_reg[29][7] ), .A1 (n_4_0_61), .A2 (n_4_0_8));
NOR2_X1 i_4_0_996 (.ZN (\partial_reg[29][6] ), .A1 (n_4_0_61), .A2 (n_4_0_7));
NOR2_X1 i_4_0_995 (.ZN (\partial_reg[29][5] ), .A1 (n_4_0_61), .A2 (n_4_0_6));
NOR2_X1 i_4_0_994 (.ZN (\partial_reg[29][4] ), .A1 (n_4_0_61), .A2 (n_4_0_5));
NOR2_X1 i_4_0_993 (.ZN (\partial_reg[29][3] ), .A1 (n_4_0_61), .A2 (n_4_0_4));
NOR2_X1 i_4_0_992 (.ZN (\partial_reg[29][2] ), .A1 (n_4_0_61), .A2 (n_4_0_3));
NOR2_X1 i_4_0_991 (.ZN (\partial_reg[29][1] ), .A1 (n_4_0_61), .A2 (n_4_0_2));
NOR2_X1 i_4_0_990 (.ZN (\partial_reg[29][0] ), .A1 (n_4_0_61), .A2 (n_4_0_1));
INV_X2 i_4_0_989 (.ZN (n_4_0_61), .A (\op2[29] ));
NOR2_X1 i_4_0_988 (.ZN (\partial_reg[28][31] ), .A1 (n_4_0_60), .A2 (n_4_0_32));
NOR2_X1 i_4_0_987 (.ZN (\partial_reg[28][30] ), .A1 (n_4_0_60), .A2 (n_4_0_31));
NOR2_X1 i_4_0_986 (.ZN (\partial_reg[28][29] ), .A1 (n_4_0_60), .A2 (n_4_0_30));
NOR2_X1 i_4_0_985 (.ZN (\partial_reg[28][28] ), .A1 (n_4_0_60), .A2 (n_4_0_29));
NOR2_X1 i_4_0_984 (.ZN (\partial_reg[28][27] ), .A1 (n_4_0_60), .A2 (n_4_0_28));
NOR2_X1 i_4_0_983 (.ZN (\partial_reg[28][26] ), .A1 (n_4_0_60), .A2 (n_4_0_27));
NOR2_X1 i_4_0_982 (.ZN (\partial_reg[28][25] ), .A1 (n_4_0_60), .A2 (n_4_0_26));
NOR2_X1 i_4_0_981 (.ZN (\partial_reg[28][24] ), .A1 (n_4_0_60), .A2 (n_4_0_25));
NOR2_X1 i_4_0_980 (.ZN (\partial_reg[28][23] ), .A1 (n_4_0_60), .A2 (n_4_0_24));
NOR2_X1 i_4_0_979 (.ZN (\partial_reg[28][22] ), .A1 (n_4_0_60), .A2 (n_4_0_23));
NOR2_X1 i_4_0_978 (.ZN (\partial_reg[28][21] ), .A1 (n_4_0_60), .A2 (n_4_0_22));
NOR2_X1 i_4_0_977 (.ZN (\partial_reg[28][20] ), .A1 (n_4_0_60), .A2 (n_4_0_21));
NOR2_X1 i_4_0_976 (.ZN (\partial_reg[28][19] ), .A1 (n_4_0_60), .A2 (n_4_0_20));
NOR2_X1 i_4_0_975 (.ZN (\partial_reg[28][18] ), .A1 (n_4_0_60), .A2 (n_4_0_19));
NOR2_X1 i_4_0_974 (.ZN (\partial_reg[28][17] ), .A1 (n_4_0_60), .A2 (n_4_0_18));
NOR2_X1 i_4_0_973 (.ZN (\partial_reg[28][16] ), .A1 (n_4_0_60), .A2 (n_4_0_17));
NOR2_X1 i_4_0_972 (.ZN (\partial_reg[28][15] ), .A1 (n_4_0_60), .A2 (n_4_0_16));
NOR2_X1 i_4_0_971 (.ZN (\partial_reg[28][14] ), .A1 (n_4_0_60), .A2 (n_4_0_15));
NOR2_X1 i_4_0_970 (.ZN (\partial_reg[28][13] ), .A1 (n_4_0_60), .A2 (n_4_0_14));
NOR2_X1 i_4_0_969 (.ZN (\partial_reg[28][12] ), .A1 (n_4_0_60), .A2 (n_4_0_13));
NOR2_X1 i_4_0_968 (.ZN (\partial_reg[28][11] ), .A1 (n_4_0_60), .A2 (n_4_0_12));
NOR2_X1 i_4_0_967 (.ZN (\partial_reg[28][10] ), .A1 (n_4_0_60), .A2 (n_4_0_11));
NOR2_X1 i_4_0_966 (.ZN (\partial_reg[28][9] ), .A1 (n_4_0_60), .A2 (n_4_0_10));
NOR2_X1 i_4_0_965 (.ZN (\partial_reg[28][8] ), .A1 (n_4_0_60), .A2 (n_4_0_9));
NOR2_X1 i_4_0_964 (.ZN (\partial_reg[28][7] ), .A1 (n_4_0_60), .A2 (n_4_0_8));
NOR2_X1 i_4_0_963 (.ZN (\partial_reg[28][6] ), .A1 (n_4_0_60), .A2 (n_4_0_7));
NOR2_X1 i_4_0_962 (.ZN (\partial_reg[28][5] ), .A1 (n_4_0_60), .A2 (n_4_0_6));
NOR2_X1 i_4_0_961 (.ZN (\partial_reg[28][4] ), .A1 (n_4_0_60), .A2 (n_4_0_5));
NOR2_X1 i_4_0_960 (.ZN (\partial_reg[28][3] ), .A1 (n_4_0_60), .A2 (n_4_0_4));
NOR2_X1 i_4_0_959 (.ZN (\partial_reg[28][2] ), .A1 (n_4_0_60), .A2 (n_4_0_3));
NOR2_X1 i_4_0_958 (.ZN (\partial_reg[28][1] ), .A1 (n_4_0_60), .A2 (n_4_0_2));
NOR2_X1 i_4_0_957 (.ZN (\partial_reg[28][0] ), .A1 (n_4_0_60), .A2 (n_4_0_1));
INV_X2 i_4_0_956 (.ZN (n_4_0_60), .A (\op2[28] ));
NOR2_X1 i_4_0_955 (.ZN (\partial_reg[27][31] ), .A1 (n_4_0_59), .A2 (n_4_0_32));
NOR2_X1 i_4_0_954 (.ZN (\partial_reg[27][30] ), .A1 (n_4_0_59), .A2 (n_4_0_31));
NOR2_X1 i_4_0_953 (.ZN (\partial_reg[27][29] ), .A1 (n_4_0_59), .A2 (n_4_0_30));
NOR2_X1 i_4_0_952 (.ZN (\partial_reg[27][28] ), .A1 (n_4_0_59), .A2 (n_4_0_29));
NOR2_X1 i_4_0_951 (.ZN (\partial_reg[27][27] ), .A1 (n_4_0_59), .A2 (n_4_0_28));
NOR2_X1 i_4_0_950 (.ZN (\partial_reg[27][26] ), .A1 (n_4_0_59), .A2 (n_4_0_27));
NOR2_X1 i_4_0_949 (.ZN (\partial_reg[27][25] ), .A1 (n_4_0_59), .A2 (n_4_0_26));
NOR2_X1 i_4_0_948 (.ZN (\partial_reg[27][24] ), .A1 (n_4_0_59), .A2 (n_4_0_25));
NOR2_X1 i_4_0_947 (.ZN (\partial_reg[27][23] ), .A1 (n_4_0_59), .A2 (n_4_0_24));
NOR2_X1 i_4_0_946 (.ZN (\partial_reg[27][22] ), .A1 (n_4_0_59), .A2 (n_4_0_23));
NOR2_X1 i_4_0_945 (.ZN (\partial_reg[27][21] ), .A1 (n_4_0_59), .A2 (n_4_0_22));
NOR2_X1 i_4_0_944 (.ZN (\partial_reg[27][20] ), .A1 (n_4_0_59), .A2 (n_4_0_21));
NOR2_X1 i_4_0_943 (.ZN (\partial_reg[27][19] ), .A1 (n_4_0_59), .A2 (n_4_0_20));
NOR2_X1 i_4_0_942 (.ZN (\partial_reg[27][18] ), .A1 (n_4_0_59), .A2 (n_4_0_19));
NOR2_X1 i_4_0_941 (.ZN (\partial_reg[27][17] ), .A1 (n_4_0_59), .A2 (n_4_0_18));
NOR2_X1 i_4_0_940 (.ZN (\partial_reg[27][16] ), .A1 (n_4_0_59), .A2 (n_4_0_17));
NOR2_X1 i_4_0_939 (.ZN (\partial_reg[27][15] ), .A1 (n_4_0_59), .A2 (n_4_0_16));
NOR2_X1 i_4_0_938 (.ZN (\partial_reg[27][14] ), .A1 (n_4_0_59), .A2 (n_4_0_15));
NOR2_X1 i_4_0_937 (.ZN (\partial_reg[27][13] ), .A1 (n_4_0_59), .A2 (n_4_0_14));
NOR2_X1 i_4_0_936 (.ZN (\partial_reg[27][12] ), .A1 (n_4_0_59), .A2 (n_4_0_13));
NOR2_X1 i_4_0_935 (.ZN (\partial_reg[27][11] ), .A1 (n_4_0_59), .A2 (n_4_0_12));
NOR2_X1 i_4_0_934 (.ZN (\partial_reg[27][10] ), .A1 (n_4_0_59), .A2 (n_4_0_11));
NOR2_X1 i_4_0_933 (.ZN (\partial_reg[27][9] ), .A1 (n_4_0_59), .A2 (n_4_0_10));
NOR2_X1 i_4_0_932 (.ZN (\partial_reg[27][8] ), .A1 (n_4_0_59), .A2 (n_4_0_9));
NOR2_X1 i_4_0_931 (.ZN (\partial_reg[27][7] ), .A1 (n_4_0_59), .A2 (n_4_0_8));
NOR2_X1 i_4_0_930 (.ZN (\partial_reg[27][6] ), .A1 (n_4_0_59), .A2 (n_4_0_7));
NOR2_X1 i_4_0_929 (.ZN (\partial_reg[27][5] ), .A1 (n_4_0_59), .A2 (n_4_0_6));
NOR2_X1 i_4_0_928 (.ZN (\partial_reg[27][4] ), .A1 (n_4_0_59), .A2 (n_4_0_5));
NOR2_X1 i_4_0_927 (.ZN (\partial_reg[27][3] ), .A1 (n_4_0_59), .A2 (n_4_0_4));
NOR2_X1 i_4_0_926 (.ZN (\partial_reg[27][2] ), .A1 (n_4_0_59), .A2 (n_4_0_3));
NOR2_X1 i_4_0_925 (.ZN (\partial_reg[27][1] ), .A1 (n_4_0_59), .A2 (n_4_0_2));
NOR2_X1 i_4_0_924 (.ZN (\partial_reg[27][0] ), .A1 (n_4_0_59), .A2 (n_4_0_1));
INV_X2 i_4_0_923 (.ZN (n_4_0_59), .A (\op2[27] ));
NOR2_X1 i_4_0_922 (.ZN (\partial_reg[26][31] ), .A1 (n_4_0_58), .A2 (n_4_0_32));
NOR2_X1 i_4_0_921 (.ZN (\partial_reg[26][30] ), .A1 (n_4_0_58), .A2 (n_4_0_31));
NOR2_X1 i_4_0_920 (.ZN (\partial_reg[26][29] ), .A1 (n_4_0_58), .A2 (n_4_0_30));
NOR2_X1 i_4_0_919 (.ZN (\partial_reg[26][28] ), .A1 (n_4_0_58), .A2 (n_4_0_29));
NOR2_X1 i_4_0_918 (.ZN (\partial_reg[26][27] ), .A1 (n_4_0_58), .A2 (n_4_0_28));
NOR2_X1 i_4_0_917 (.ZN (\partial_reg[26][26] ), .A1 (n_4_0_58), .A2 (n_4_0_27));
NOR2_X1 i_4_0_916 (.ZN (\partial_reg[26][25] ), .A1 (n_4_0_58), .A2 (n_4_0_26));
NOR2_X1 i_4_0_915 (.ZN (\partial_reg[26][24] ), .A1 (n_4_0_58), .A2 (n_4_0_25));
NOR2_X1 i_4_0_914 (.ZN (\partial_reg[26][23] ), .A1 (n_4_0_58), .A2 (n_4_0_24));
NOR2_X1 i_4_0_913 (.ZN (\partial_reg[26][22] ), .A1 (n_4_0_58), .A2 (n_4_0_23));
NOR2_X1 i_4_0_912 (.ZN (\partial_reg[26][21] ), .A1 (n_4_0_58), .A2 (n_4_0_22));
NOR2_X1 i_4_0_911 (.ZN (\partial_reg[26][20] ), .A1 (n_4_0_58), .A2 (n_4_0_21));
NOR2_X1 i_4_0_910 (.ZN (\partial_reg[26][19] ), .A1 (n_4_0_58), .A2 (n_4_0_20));
NOR2_X1 i_4_0_909 (.ZN (\partial_reg[26][18] ), .A1 (n_4_0_58), .A2 (n_4_0_19));
NOR2_X1 i_4_0_908 (.ZN (\partial_reg[26][17] ), .A1 (n_4_0_58), .A2 (n_4_0_18));
NOR2_X1 i_4_0_907 (.ZN (\partial_reg[26][16] ), .A1 (n_4_0_58), .A2 (n_4_0_17));
NOR2_X1 i_4_0_906 (.ZN (\partial_reg[26][15] ), .A1 (n_4_0_58), .A2 (n_4_0_16));
NOR2_X1 i_4_0_905 (.ZN (\partial_reg[26][14] ), .A1 (n_4_0_58), .A2 (n_4_0_15));
NOR2_X1 i_4_0_904 (.ZN (\partial_reg[26][13] ), .A1 (n_4_0_58), .A2 (n_4_0_14));
NOR2_X1 i_4_0_903 (.ZN (\partial_reg[26][12] ), .A1 (n_4_0_58), .A2 (n_4_0_13));
NOR2_X1 i_4_0_902 (.ZN (\partial_reg[26][11] ), .A1 (n_4_0_58), .A2 (n_4_0_12));
NOR2_X1 i_4_0_901 (.ZN (\partial_reg[26][10] ), .A1 (n_4_0_58), .A2 (n_4_0_11));
NOR2_X1 i_4_0_900 (.ZN (\partial_reg[26][9] ), .A1 (n_4_0_58), .A2 (n_4_0_10));
NOR2_X1 i_4_0_899 (.ZN (\partial_reg[26][8] ), .A1 (n_4_0_58), .A2 (n_4_0_9));
NOR2_X1 i_4_0_898 (.ZN (\partial_reg[26][7] ), .A1 (n_4_0_58), .A2 (n_4_0_8));
NOR2_X1 i_4_0_897 (.ZN (\partial_reg[26][6] ), .A1 (n_4_0_58), .A2 (n_4_0_7));
NOR2_X1 i_4_0_896 (.ZN (\partial_reg[26][5] ), .A1 (n_4_0_58), .A2 (n_4_0_6));
NOR2_X1 i_4_0_895 (.ZN (\partial_reg[26][4] ), .A1 (n_4_0_58), .A2 (n_4_0_5));
NOR2_X1 i_4_0_894 (.ZN (\partial_reg[26][3] ), .A1 (n_4_0_58), .A2 (n_4_0_4));
NOR2_X1 i_4_0_893 (.ZN (\partial_reg[26][2] ), .A1 (n_4_0_58), .A2 (n_4_0_3));
NOR2_X1 i_4_0_892 (.ZN (\partial_reg[26][1] ), .A1 (n_4_0_58), .A2 (n_4_0_2));
NOR2_X1 i_4_0_891 (.ZN (\partial_reg[26][0] ), .A1 (n_4_0_58), .A2 (n_4_0_1));
INV_X2 i_4_0_890 (.ZN (n_4_0_58), .A (\op2[26] ));
NOR2_X1 i_4_0_889 (.ZN (\partial_reg[25][31] ), .A1 (n_4_0_57), .A2 (n_4_0_32));
NOR2_X1 i_4_0_888 (.ZN (\partial_reg[25][30] ), .A1 (n_4_0_57), .A2 (n_4_0_31));
NOR2_X1 i_4_0_887 (.ZN (\partial_reg[25][29] ), .A1 (n_4_0_57), .A2 (n_4_0_30));
NOR2_X1 i_4_0_886 (.ZN (\partial_reg[25][28] ), .A1 (n_4_0_57), .A2 (n_4_0_29));
NOR2_X1 i_4_0_885 (.ZN (\partial_reg[25][27] ), .A1 (n_4_0_57), .A2 (n_4_0_28));
NOR2_X1 i_4_0_884 (.ZN (\partial_reg[25][26] ), .A1 (n_4_0_57), .A2 (n_4_0_27));
NOR2_X1 i_4_0_883 (.ZN (\partial_reg[25][25] ), .A1 (n_4_0_57), .A2 (n_4_0_26));
NOR2_X1 i_4_0_882 (.ZN (\partial_reg[25][24] ), .A1 (n_4_0_57), .A2 (n_4_0_25));
NOR2_X1 i_4_0_881 (.ZN (\partial_reg[25][23] ), .A1 (n_4_0_57), .A2 (n_4_0_24));
NOR2_X1 i_4_0_880 (.ZN (\partial_reg[25][22] ), .A1 (n_4_0_57), .A2 (n_4_0_23));
NOR2_X1 i_4_0_879 (.ZN (\partial_reg[25][21] ), .A1 (n_4_0_57), .A2 (n_4_0_22));
NOR2_X1 i_4_0_878 (.ZN (\partial_reg[25][20] ), .A1 (n_4_0_57), .A2 (n_4_0_21));
NOR2_X1 i_4_0_877 (.ZN (\partial_reg[25][19] ), .A1 (n_4_0_57), .A2 (n_4_0_20));
NOR2_X1 i_4_0_876 (.ZN (\partial_reg[25][18] ), .A1 (n_4_0_57), .A2 (n_4_0_19));
NOR2_X1 i_4_0_875 (.ZN (\partial_reg[25][17] ), .A1 (n_4_0_57), .A2 (n_4_0_18));
NOR2_X1 i_4_0_874 (.ZN (\partial_reg[25][16] ), .A1 (n_4_0_57), .A2 (n_4_0_17));
NOR2_X1 i_4_0_873 (.ZN (\partial_reg[25][15] ), .A1 (n_4_0_57), .A2 (n_4_0_16));
NOR2_X1 i_4_0_872 (.ZN (\partial_reg[25][14] ), .A1 (n_4_0_57), .A2 (n_4_0_15));
NOR2_X1 i_4_0_871 (.ZN (\partial_reg[25][13] ), .A1 (n_4_0_57), .A2 (n_4_0_14));
NOR2_X1 i_4_0_870 (.ZN (\partial_reg[25][12] ), .A1 (n_4_0_57), .A2 (n_4_0_13));
NOR2_X1 i_4_0_869 (.ZN (\partial_reg[25][11] ), .A1 (n_4_0_57), .A2 (n_4_0_12));
NOR2_X1 i_4_0_868 (.ZN (\partial_reg[25][10] ), .A1 (n_4_0_57), .A2 (n_4_0_11));
NOR2_X1 i_4_0_867 (.ZN (\partial_reg[25][9] ), .A1 (n_4_0_57), .A2 (n_4_0_10));
NOR2_X1 i_4_0_866 (.ZN (\partial_reg[25][8] ), .A1 (n_4_0_57), .A2 (n_4_0_9));
NOR2_X1 i_4_0_865 (.ZN (\partial_reg[25][7] ), .A1 (n_4_0_57), .A2 (n_4_0_8));
NOR2_X1 i_4_0_864 (.ZN (\partial_reg[25][6] ), .A1 (n_4_0_57), .A2 (n_4_0_7));
NOR2_X1 i_4_0_863 (.ZN (\partial_reg[25][5] ), .A1 (n_4_0_57), .A2 (n_4_0_6));
NOR2_X1 i_4_0_862 (.ZN (\partial_reg[25][4] ), .A1 (n_4_0_57), .A2 (n_4_0_5));
NOR2_X1 i_4_0_861 (.ZN (\partial_reg[25][3] ), .A1 (n_4_0_57), .A2 (n_4_0_4));
NOR2_X1 i_4_0_860 (.ZN (\partial_reg[25][2] ), .A1 (n_4_0_57), .A2 (n_4_0_3));
NOR2_X1 i_4_0_859 (.ZN (\partial_reg[25][1] ), .A1 (n_4_0_57), .A2 (n_4_0_2));
NOR2_X1 i_4_0_858 (.ZN (\partial_reg[25][0] ), .A1 (n_4_0_57), .A2 (n_4_0_1));
INV_X2 i_4_0_857 (.ZN (n_4_0_57), .A (\op2[25] ));
NOR2_X1 i_4_0_856 (.ZN (\partial_reg[24][31] ), .A1 (n_4_0_56), .A2 (n_4_0_32));
NOR2_X1 i_4_0_855 (.ZN (\partial_reg[24][30] ), .A1 (n_4_0_56), .A2 (n_4_0_31));
NOR2_X1 i_4_0_854 (.ZN (\partial_reg[24][29] ), .A1 (n_4_0_56), .A2 (n_4_0_30));
NOR2_X1 i_4_0_853 (.ZN (\partial_reg[24][28] ), .A1 (n_4_0_56), .A2 (n_4_0_29));
NOR2_X1 i_4_0_852 (.ZN (\partial_reg[24][27] ), .A1 (n_4_0_56), .A2 (n_4_0_28));
NOR2_X1 i_4_0_851 (.ZN (\partial_reg[24][26] ), .A1 (n_4_0_56), .A2 (n_4_0_27));
NOR2_X1 i_4_0_850 (.ZN (\partial_reg[24][25] ), .A1 (n_4_0_56), .A2 (n_4_0_26));
NOR2_X1 i_4_0_849 (.ZN (\partial_reg[24][24] ), .A1 (n_4_0_56), .A2 (n_4_0_25));
NOR2_X1 i_4_0_848 (.ZN (\partial_reg[24][23] ), .A1 (n_4_0_56), .A2 (n_4_0_24));
NOR2_X1 i_4_0_847 (.ZN (\partial_reg[24][22] ), .A1 (n_4_0_56), .A2 (n_4_0_23));
NOR2_X1 i_4_0_846 (.ZN (\partial_reg[24][21] ), .A1 (n_4_0_56), .A2 (n_4_0_22));
NOR2_X1 i_4_0_845 (.ZN (\partial_reg[24][20] ), .A1 (n_4_0_56), .A2 (n_4_0_21));
NOR2_X1 i_4_0_844 (.ZN (\partial_reg[24][19] ), .A1 (n_4_0_56), .A2 (n_4_0_20));
NOR2_X1 i_4_0_843 (.ZN (\partial_reg[24][18] ), .A1 (n_4_0_56), .A2 (n_4_0_19));
NOR2_X1 i_4_0_842 (.ZN (\partial_reg[24][17] ), .A1 (n_4_0_56), .A2 (n_4_0_18));
NOR2_X1 i_4_0_841 (.ZN (\partial_reg[24][16] ), .A1 (n_4_0_56), .A2 (n_4_0_17));
NOR2_X1 i_4_0_840 (.ZN (\partial_reg[24][15] ), .A1 (n_4_0_56), .A2 (n_4_0_16));
NOR2_X1 i_4_0_839 (.ZN (\partial_reg[24][14] ), .A1 (n_4_0_56), .A2 (n_4_0_15));
NOR2_X1 i_4_0_838 (.ZN (\partial_reg[24][13] ), .A1 (n_4_0_56), .A2 (n_4_0_14));
NOR2_X1 i_4_0_837 (.ZN (\partial_reg[24][12] ), .A1 (n_4_0_56), .A2 (n_4_0_13));
NOR2_X1 i_4_0_836 (.ZN (\partial_reg[24][11] ), .A1 (n_4_0_56), .A2 (n_4_0_12));
NOR2_X1 i_4_0_835 (.ZN (\partial_reg[24][10] ), .A1 (n_4_0_56), .A2 (n_4_0_11));
NOR2_X1 i_4_0_834 (.ZN (\partial_reg[24][9] ), .A1 (n_4_0_56), .A2 (n_4_0_10));
NOR2_X1 i_4_0_833 (.ZN (\partial_reg[24][8] ), .A1 (n_4_0_56), .A2 (n_4_0_9));
NOR2_X1 i_4_0_832 (.ZN (\partial_reg[24][7] ), .A1 (n_4_0_56), .A2 (n_4_0_8));
NOR2_X1 i_4_0_831 (.ZN (\partial_reg[24][6] ), .A1 (n_4_0_56), .A2 (n_4_0_7));
NOR2_X1 i_4_0_830 (.ZN (\partial_reg[24][5] ), .A1 (n_4_0_56), .A2 (n_4_0_6));
NOR2_X1 i_4_0_829 (.ZN (\partial_reg[24][4] ), .A1 (n_4_0_56), .A2 (n_4_0_5));
NOR2_X1 i_4_0_828 (.ZN (\partial_reg[24][3] ), .A1 (n_4_0_56), .A2 (n_4_0_4));
NOR2_X1 i_4_0_827 (.ZN (\partial_reg[24][2] ), .A1 (n_4_0_56), .A2 (n_4_0_3));
NOR2_X1 i_4_0_826 (.ZN (\partial_reg[24][1] ), .A1 (n_4_0_56), .A2 (n_4_0_2));
NOR2_X1 i_4_0_825 (.ZN (\partial_reg[24][0] ), .A1 (n_4_0_56), .A2 (n_4_0_1));
INV_X2 i_4_0_824 (.ZN (n_4_0_56), .A (\op2[24] ));
NOR2_X1 i_4_0_823 (.ZN (\partial_reg[23][31] ), .A1 (n_4_0_55), .A2 (n_4_0_32));
NOR2_X1 i_4_0_822 (.ZN (\partial_reg[23][30] ), .A1 (n_4_0_55), .A2 (n_4_0_31));
NOR2_X1 i_4_0_821 (.ZN (\partial_reg[23][29] ), .A1 (n_4_0_55), .A2 (n_4_0_30));
NOR2_X1 i_4_0_820 (.ZN (\partial_reg[23][28] ), .A1 (n_4_0_55), .A2 (n_4_0_29));
NOR2_X1 i_4_0_819 (.ZN (\partial_reg[23][27] ), .A1 (n_4_0_55), .A2 (n_4_0_28));
NOR2_X1 i_4_0_818 (.ZN (\partial_reg[23][26] ), .A1 (n_4_0_55), .A2 (n_4_0_27));
NOR2_X1 i_4_0_817 (.ZN (\partial_reg[23][25] ), .A1 (n_4_0_55), .A2 (n_4_0_26));
NOR2_X1 i_4_0_816 (.ZN (\partial_reg[23][24] ), .A1 (n_4_0_55), .A2 (n_4_0_25));
NOR2_X1 i_4_0_815 (.ZN (\partial_reg[23][23] ), .A1 (n_4_0_55), .A2 (n_4_0_24));
NOR2_X1 i_4_0_814 (.ZN (\partial_reg[23][22] ), .A1 (n_4_0_55), .A2 (n_4_0_23));
NOR2_X1 i_4_0_813 (.ZN (\partial_reg[23][21] ), .A1 (n_4_0_55), .A2 (n_4_0_22));
NOR2_X1 i_4_0_812 (.ZN (\partial_reg[23][20] ), .A1 (n_4_0_55), .A2 (n_4_0_21));
NOR2_X1 i_4_0_811 (.ZN (\partial_reg[23][19] ), .A1 (n_4_0_55), .A2 (n_4_0_20));
NOR2_X1 i_4_0_810 (.ZN (\partial_reg[23][18] ), .A1 (n_4_0_55), .A2 (n_4_0_19));
NOR2_X1 i_4_0_809 (.ZN (\partial_reg[23][17] ), .A1 (n_4_0_55), .A2 (n_4_0_18));
NOR2_X1 i_4_0_808 (.ZN (\partial_reg[23][16] ), .A1 (n_4_0_55), .A2 (n_4_0_17));
NOR2_X1 i_4_0_807 (.ZN (\partial_reg[23][15] ), .A1 (n_4_0_55), .A2 (n_4_0_16));
NOR2_X1 i_4_0_806 (.ZN (\partial_reg[23][14] ), .A1 (n_4_0_55), .A2 (n_4_0_15));
NOR2_X1 i_4_0_805 (.ZN (\partial_reg[23][13] ), .A1 (n_4_0_55), .A2 (n_4_0_14));
NOR2_X1 i_4_0_804 (.ZN (\partial_reg[23][12] ), .A1 (n_4_0_55), .A2 (n_4_0_13));
NOR2_X1 i_4_0_803 (.ZN (\partial_reg[23][11] ), .A1 (n_4_0_55), .A2 (n_4_0_12));
NOR2_X1 i_4_0_802 (.ZN (\partial_reg[23][10] ), .A1 (n_4_0_55), .A2 (n_4_0_11));
NOR2_X1 i_4_0_801 (.ZN (\partial_reg[23][9] ), .A1 (n_4_0_55), .A2 (n_4_0_10));
NOR2_X1 i_4_0_800 (.ZN (\partial_reg[23][8] ), .A1 (n_4_0_55), .A2 (n_4_0_9));
NOR2_X1 i_4_0_799 (.ZN (\partial_reg[23][7] ), .A1 (n_4_0_55), .A2 (n_4_0_8));
NOR2_X1 i_4_0_798 (.ZN (\partial_reg[23][6] ), .A1 (n_4_0_55), .A2 (n_4_0_7));
NOR2_X1 i_4_0_797 (.ZN (\partial_reg[23][5] ), .A1 (n_4_0_55), .A2 (n_4_0_6));
NOR2_X1 i_4_0_796 (.ZN (\partial_reg[23][4] ), .A1 (n_4_0_55), .A2 (n_4_0_5));
NOR2_X1 i_4_0_795 (.ZN (\partial_reg[23][3] ), .A1 (n_4_0_55), .A2 (n_4_0_4));
NOR2_X1 i_4_0_794 (.ZN (\partial_reg[23][2] ), .A1 (n_4_0_55), .A2 (n_4_0_3));
NOR2_X1 i_4_0_793 (.ZN (\partial_reg[23][1] ), .A1 (n_4_0_55), .A2 (n_4_0_2));
NOR2_X1 i_4_0_792 (.ZN (\partial_reg[23][0] ), .A1 (n_4_0_55), .A2 (n_4_0_1));
INV_X2 i_4_0_791 (.ZN (n_4_0_55), .A (\op2[23] ));
NOR2_X1 i_4_0_790 (.ZN (\partial_reg[22][31] ), .A1 (n_4_0_54), .A2 (n_4_0_32));
NOR2_X1 i_4_0_789 (.ZN (\partial_reg[22][30] ), .A1 (n_4_0_54), .A2 (n_4_0_31));
NOR2_X1 i_4_0_788 (.ZN (\partial_reg[22][29] ), .A1 (n_4_0_54), .A2 (n_4_0_30));
NOR2_X1 i_4_0_787 (.ZN (\partial_reg[22][28] ), .A1 (n_4_0_54), .A2 (n_4_0_29));
NOR2_X1 i_4_0_786 (.ZN (\partial_reg[22][27] ), .A1 (n_4_0_54), .A2 (n_4_0_28));
NOR2_X1 i_4_0_785 (.ZN (\partial_reg[22][26] ), .A1 (n_4_0_54), .A2 (n_4_0_27));
NOR2_X1 i_4_0_784 (.ZN (\partial_reg[22][25] ), .A1 (n_4_0_54), .A2 (n_4_0_26));
NOR2_X1 i_4_0_783 (.ZN (\partial_reg[22][24] ), .A1 (n_4_0_54), .A2 (n_4_0_25));
NOR2_X1 i_4_0_782 (.ZN (\partial_reg[22][23] ), .A1 (n_4_0_54), .A2 (n_4_0_24));
NOR2_X1 i_4_0_781 (.ZN (\partial_reg[22][22] ), .A1 (n_4_0_54), .A2 (n_4_0_23));
NOR2_X1 i_4_0_780 (.ZN (\partial_reg[22][21] ), .A1 (n_4_0_54), .A2 (n_4_0_22));
NOR2_X1 i_4_0_779 (.ZN (\partial_reg[22][20] ), .A1 (n_4_0_54), .A2 (n_4_0_21));
NOR2_X1 i_4_0_778 (.ZN (\partial_reg[22][19] ), .A1 (n_4_0_54), .A2 (n_4_0_20));
NOR2_X1 i_4_0_777 (.ZN (\partial_reg[22][18] ), .A1 (n_4_0_54), .A2 (n_4_0_19));
NOR2_X1 i_4_0_776 (.ZN (\partial_reg[22][17] ), .A1 (n_4_0_54), .A2 (n_4_0_18));
NOR2_X1 i_4_0_775 (.ZN (\partial_reg[22][16] ), .A1 (n_4_0_54), .A2 (n_4_0_17));
NOR2_X1 i_4_0_774 (.ZN (\partial_reg[22][15] ), .A1 (n_4_0_54), .A2 (n_4_0_16));
NOR2_X1 i_4_0_773 (.ZN (\partial_reg[22][14] ), .A1 (n_4_0_54), .A2 (n_4_0_15));
NOR2_X1 i_4_0_772 (.ZN (\partial_reg[22][13] ), .A1 (n_4_0_54), .A2 (n_4_0_14));
NOR2_X1 i_4_0_771 (.ZN (\partial_reg[22][12] ), .A1 (n_4_0_54), .A2 (n_4_0_13));
NOR2_X1 i_4_0_770 (.ZN (\partial_reg[22][11] ), .A1 (n_4_0_54), .A2 (n_4_0_12));
NOR2_X1 i_4_0_769 (.ZN (\partial_reg[22][10] ), .A1 (n_4_0_54), .A2 (n_4_0_11));
NOR2_X1 i_4_0_768 (.ZN (\partial_reg[22][9] ), .A1 (n_4_0_54), .A2 (n_4_0_10));
NOR2_X1 i_4_0_767 (.ZN (\partial_reg[22][8] ), .A1 (n_4_0_54), .A2 (n_4_0_9));
NOR2_X1 i_4_0_766 (.ZN (\partial_reg[22][7] ), .A1 (n_4_0_54), .A2 (n_4_0_8));
NOR2_X1 i_4_0_765 (.ZN (\partial_reg[22][6] ), .A1 (n_4_0_54), .A2 (n_4_0_7));
NOR2_X1 i_4_0_764 (.ZN (\partial_reg[22][5] ), .A1 (n_4_0_54), .A2 (n_4_0_6));
NOR2_X1 i_4_0_763 (.ZN (\partial_reg[22][4] ), .A1 (n_4_0_54), .A2 (n_4_0_5));
NOR2_X1 i_4_0_762 (.ZN (\partial_reg[22][3] ), .A1 (n_4_0_54), .A2 (n_4_0_4));
NOR2_X1 i_4_0_761 (.ZN (\partial_reg[22][2] ), .A1 (n_4_0_54), .A2 (n_4_0_3));
NOR2_X1 i_4_0_760 (.ZN (\partial_reg[22][1] ), .A1 (n_4_0_54), .A2 (n_4_0_2));
NOR2_X1 i_4_0_759 (.ZN (\partial_reg[22][0] ), .A1 (n_4_0_54), .A2 (n_4_0_1));
INV_X2 i_4_0_758 (.ZN (n_4_0_54), .A (\op2[22] ));
NOR2_X1 i_4_0_757 (.ZN (\partial_reg[21][31] ), .A1 (n_4_0_53), .A2 (n_4_0_32));
NOR2_X1 i_4_0_756 (.ZN (\partial_reg[21][30] ), .A1 (n_4_0_53), .A2 (n_4_0_31));
NOR2_X1 i_4_0_755 (.ZN (\partial_reg[21][29] ), .A1 (n_4_0_53), .A2 (n_4_0_30));
NOR2_X1 i_4_0_754 (.ZN (\partial_reg[21][28] ), .A1 (n_4_0_53), .A2 (n_4_0_29));
NOR2_X1 i_4_0_753 (.ZN (\partial_reg[21][27] ), .A1 (n_4_0_53), .A2 (n_4_0_28));
NOR2_X1 i_4_0_752 (.ZN (\partial_reg[21][26] ), .A1 (n_4_0_53), .A2 (n_4_0_27));
NOR2_X1 i_4_0_751 (.ZN (\partial_reg[21][25] ), .A1 (n_4_0_53), .A2 (n_4_0_26));
NOR2_X1 i_4_0_750 (.ZN (\partial_reg[21][24] ), .A1 (n_4_0_53), .A2 (n_4_0_25));
NOR2_X1 i_4_0_749 (.ZN (\partial_reg[21][23] ), .A1 (n_4_0_53), .A2 (n_4_0_24));
NOR2_X1 i_4_0_748 (.ZN (\partial_reg[21][22] ), .A1 (n_4_0_53), .A2 (n_4_0_23));
NOR2_X1 i_4_0_747 (.ZN (\partial_reg[21][21] ), .A1 (n_4_0_53), .A2 (n_4_0_22));
NOR2_X1 i_4_0_746 (.ZN (\partial_reg[21][20] ), .A1 (n_4_0_53), .A2 (n_4_0_21));
NOR2_X1 i_4_0_745 (.ZN (\partial_reg[21][19] ), .A1 (n_4_0_53), .A2 (n_4_0_20));
NOR2_X1 i_4_0_744 (.ZN (\partial_reg[21][18] ), .A1 (n_4_0_53), .A2 (n_4_0_19));
NOR2_X1 i_4_0_743 (.ZN (\partial_reg[21][17] ), .A1 (n_4_0_53), .A2 (n_4_0_18));
NOR2_X1 i_4_0_742 (.ZN (\partial_reg[21][16] ), .A1 (n_4_0_53), .A2 (n_4_0_17));
NOR2_X1 i_4_0_741 (.ZN (\partial_reg[21][15] ), .A1 (n_4_0_53), .A2 (n_4_0_16));
NOR2_X1 i_4_0_740 (.ZN (\partial_reg[21][14] ), .A1 (n_4_0_53), .A2 (n_4_0_15));
NOR2_X1 i_4_0_739 (.ZN (\partial_reg[21][13] ), .A1 (n_4_0_53), .A2 (n_4_0_14));
NOR2_X1 i_4_0_738 (.ZN (\partial_reg[21][12] ), .A1 (n_4_0_53), .A2 (n_4_0_13));
NOR2_X1 i_4_0_737 (.ZN (\partial_reg[21][11] ), .A1 (n_4_0_53), .A2 (n_4_0_12));
NOR2_X1 i_4_0_736 (.ZN (\partial_reg[21][10] ), .A1 (n_4_0_53), .A2 (n_4_0_11));
NOR2_X1 i_4_0_735 (.ZN (\partial_reg[21][9] ), .A1 (n_4_0_53), .A2 (n_4_0_10));
NOR2_X1 i_4_0_734 (.ZN (\partial_reg[21][8] ), .A1 (n_4_0_53), .A2 (n_4_0_9));
NOR2_X1 i_4_0_733 (.ZN (\partial_reg[21][7] ), .A1 (n_4_0_53), .A2 (n_4_0_8));
NOR2_X1 i_4_0_732 (.ZN (\partial_reg[21][6] ), .A1 (n_4_0_53), .A2 (n_4_0_7));
NOR2_X1 i_4_0_731 (.ZN (\partial_reg[21][5] ), .A1 (n_4_0_53), .A2 (n_4_0_6));
NOR2_X1 i_4_0_730 (.ZN (\partial_reg[21][4] ), .A1 (n_4_0_53), .A2 (n_4_0_5));
NOR2_X1 i_4_0_729 (.ZN (\partial_reg[21][3] ), .A1 (n_4_0_53), .A2 (n_4_0_4));
NOR2_X1 i_4_0_728 (.ZN (\partial_reg[21][2] ), .A1 (n_4_0_53), .A2 (n_4_0_3));
NOR2_X1 i_4_0_727 (.ZN (\partial_reg[21][1] ), .A1 (n_4_0_53), .A2 (n_4_0_2));
NOR2_X1 i_4_0_726 (.ZN (\partial_reg[21][0] ), .A1 (n_4_0_53), .A2 (n_4_0_1));
INV_X2 i_4_0_725 (.ZN (n_4_0_53), .A (\op2[21] ));
NOR2_X1 i_4_0_724 (.ZN (\partial_reg[20][31] ), .A1 (n_4_0_52), .A2 (n_4_0_32));
NOR2_X1 i_4_0_723 (.ZN (\partial_reg[20][30] ), .A1 (n_4_0_52), .A2 (n_4_0_31));
NOR2_X1 i_4_0_722 (.ZN (\partial_reg[20][29] ), .A1 (n_4_0_52), .A2 (n_4_0_30));
NOR2_X1 i_4_0_721 (.ZN (\partial_reg[20][28] ), .A1 (n_4_0_52), .A2 (n_4_0_29));
NOR2_X1 i_4_0_720 (.ZN (\partial_reg[20][27] ), .A1 (n_4_0_52), .A2 (n_4_0_28));
NOR2_X1 i_4_0_719 (.ZN (\partial_reg[20][26] ), .A1 (n_4_0_52), .A2 (n_4_0_27));
NOR2_X1 i_4_0_718 (.ZN (\partial_reg[20][25] ), .A1 (n_4_0_52), .A2 (n_4_0_26));
NOR2_X1 i_4_0_717 (.ZN (\partial_reg[20][24] ), .A1 (n_4_0_52), .A2 (n_4_0_25));
NOR2_X1 i_4_0_716 (.ZN (\partial_reg[20][23] ), .A1 (n_4_0_52), .A2 (n_4_0_24));
NOR2_X1 i_4_0_715 (.ZN (\partial_reg[20][22] ), .A1 (n_4_0_52), .A2 (n_4_0_23));
NOR2_X1 i_4_0_714 (.ZN (\partial_reg[20][21] ), .A1 (n_4_0_52), .A2 (n_4_0_22));
NOR2_X1 i_4_0_713 (.ZN (\partial_reg[20][20] ), .A1 (n_4_0_52), .A2 (n_4_0_21));
NOR2_X1 i_4_0_712 (.ZN (\partial_reg[20][19] ), .A1 (n_4_0_52), .A2 (n_4_0_20));
NOR2_X1 i_4_0_711 (.ZN (\partial_reg[20][18] ), .A1 (n_4_0_52), .A2 (n_4_0_19));
NOR2_X1 i_4_0_710 (.ZN (\partial_reg[20][17] ), .A1 (n_4_0_52), .A2 (n_4_0_18));
NOR2_X1 i_4_0_709 (.ZN (\partial_reg[20][16] ), .A1 (n_4_0_52), .A2 (n_4_0_17));
NOR2_X1 i_4_0_708 (.ZN (\partial_reg[20][15] ), .A1 (n_4_0_52), .A2 (n_4_0_16));
NOR2_X1 i_4_0_707 (.ZN (\partial_reg[20][14] ), .A1 (n_4_0_52), .A2 (n_4_0_15));
NOR2_X1 i_4_0_706 (.ZN (\partial_reg[20][13] ), .A1 (n_4_0_52), .A2 (n_4_0_14));
NOR2_X1 i_4_0_705 (.ZN (\partial_reg[20][12] ), .A1 (n_4_0_52), .A2 (n_4_0_13));
NOR2_X1 i_4_0_704 (.ZN (\partial_reg[20][11] ), .A1 (n_4_0_52), .A2 (n_4_0_12));
NOR2_X1 i_4_0_703 (.ZN (\partial_reg[20][10] ), .A1 (n_4_0_52), .A2 (n_4_0_11));
NOR2_X1 i_4_0_702 (.ZN (\partial_reg[20][9] ), .A1 (n_4_0_52), .A2 (n_4_0_10));
NOR2_X1 i_4_0_701 (.ZN (\partial_reg[20][8] ), .A1 (n_4_0_52), .A2 (n_4_0_9));
NOR2_X1 i_4_0_700 (.ZN (\partial_reg[20][7] ), .A1 (n_4_0_52), .A2 (n_4_0_8));
NOR2_X1 i_4_0_699 (.ZN (\partial_reg[20][6] ), .A1 (n_4_0_52), .A2 (n_4_0_7));
NOR2_X1 i_4_0_698 (.ZN (\partial_reg[20][5] ), .A1 (n_4_0_52), .A2 (n_4_0_6));
NOR2_X1 i_4_0_697 (.ZN (\partial_reg[20][4] ), .A1 (n_4_0_52), .A2 (n_4_0_5));
NOR2_X1 i_4_0_696 (.ZN (\partial_reg[20][3] ), .A1 (n_4_0_52), .A2 (n_4_0_4));
NOR2_X1 i_4_0_695 (.ZN (\partial_reg[20][2] ), .A1 (n_4_0_52), .A2 (n_4_0_3));
NOR2_X1 i_4_0_694 (.ZN (\partial_reg[20][1] ), .A1 (n_4_0_52), .A2 (n_4_0_2));
NOR2_X1 i_4_0_693 (.ZN (\partial_reg[20][0] ), .A1 (n_4_0_52), .A2 (n_4_0_1));
INV_X2 i_4_0_692 (.ZN (n_4_0_52), .A (\op2[20] ));
NOR2_X1 i_4_0_691 (.ZN (\partial_reg[19][31] ), .A1 (n_4_0_51), .A2 (n_4_0_32));
NOR2_X1 i_4_0_690 (.ZN (\partial_reg[19][30] ), .A1 (n_4_0_51), .A2 (n_4_0_31));
NOR2_X1 i_4_0_689 (.ZN (\partial_reg[19][29] ), .A1 (n_4_0_51), .A2 (n_4_0_30));
NOR2_X1 i_4_0_688 (.ZN (\partial_reg[19][28] ), .A1 (n_4_0_51), .A2 (n_4_0_29));
NOR2_X1 i_4_0_687 (.ZN (\partial_reg[19][27] ), .A1 (n_4_0_51), .A2 (n_4_0_28));
NOR2_X1 i_4_0_686 (.ZN (\partial_reg[19][26] ), .A1 (n_4_0_51), .A2 (n_4_0_27));
NOR2_X1 i_4_0_685 (.ZN (\partial_reg[19][25] ), .A1 (n_4_0_51), .A2 (n_4_0_26));
NOR2_X1 i_4_0_684 (.ZN (\partial_reg[19][24] ), .A1 (n_4_0_51), .A2 (n_4_0_25));
NOR2_X1 i_4_0_683 (.ZN (\partial_reg[19][23] ), .A1 (n_4_0_51), .A2 (n_4_0_24));
NOR2_X1 i_4_0_682 (.ZN (\partial_reg[19][22] ), .A1 (n_4_0_51), .A2 (n_4_0_23));
NOR2_X1 i_4_0_681 (.ZN (\partial_reg[19][21] ), .A1 (n_4_0_51), .A2 (n_4_0_22));
NOR2_X1 i_4_0_680 (.ZN (\partial_reg[19][20] ), .A1 (n_4_0_51), .A2 (n_4_0_21));
NOR2_X1 i_4_0_679 (.ZN (\partial_reg[19][19] ), .A1 (n_4_0_51), .A2 (n_4_0_20));
NOR2_X1 i_4_0_678 (.ZN (\partial_reg[19][18] ), .A1 (n_4_0_51), .A2 (n_4_0_19));
NOR2_X1 i_4_0_677 (.ZN (\partial_reg[19][17] ), .A1 (n_4_0_51), .A2 (n_4_0_18));
NOR2_X1 i_4_0_676 (.ZN (\partial_reg[19][16] ), .A1 (n_4_0_51), .A2 (n_4_0_17));
NOR2_X1 i_4_0_675 (.ZN (\partial_reg[19][15] ), .A1 (n_4_0_51), .A2 (n_4_0_16));
NOR2_X1 i_4_0_674 (.ZN (\partial_reg[19][14] ), .A1 (n_4_0_51), .A2 (n_4_0_15));
NOR2_X1 i_4_0_673 (.ZN (\partial_reg[19][13] ), .A1 (n_4_0_51), .A2 (n_4_0_14));
NOR2_X1 i_4_0_672 (.ZN (\partial_reg[19][12] ), .A1 (n_4_0_51), .A2 (n_4_0_13));
NOR2_X1 i_4_0_671 (.ZN (\partial_reg[19][11] ), .A1 (n_4_0_51), .A2 (n_4_0_12));
NOR2_X1 i_4_0_670 (.ZN (\partial_reg[19][10] ), .A1 (n_4_0_51), .A2 (n_4_0_11));
NOR2_X1 i_4_0_669 (.ZN (\partial_reg[19][9] ), .A1 (n_4_0_51), .A2 (n_4_0_10));
NOR2_X1 i_4_0_668 (.ZN (\partial_reg[19][8] ), .A1 (n_4_0_51), .A2 (n_4_0_9));
NOR2_X1 i_4_0_667 (.ZN (\partial_reg[19][7] ), .A1 (n_4_0_51), .A2 (n_4_0_8));
NOR2_X1 i_4_0_666 (.ZN (\partial_reg[19][6] ), .A1 (n_4_0_51), .A2 (n_4_0_7));
NOR2_X1 i_4_0_665 (.ZN (\partial_reg[19][5] ), .A1 (n_4_0_51), .A2 (n_4_0_6));
NOR2_X1 i_4_0_664 (.ZN (\partial_reg[19][4] ), .A1 (n_4_0_51), .A2 (n_4_0_5));
NOR2_X1 i_4_0_663 (.ZN (\partial_reg[19][3] ), .A1 (n_4_0_51), .A2 (n_4_0_4));
NOR2_X1 i_4_0_662 (.ZN (\partial_reg[19][2] ), .A1 (n_4_0_51), .A2 (n_4_0_3));
NOR2_X1 i_4_0_661 (.ZN (\partial_reg[19][1] ), .A1 (n_4_0_51), .A2 (n_4_0_2));
NOR2_X1 i_4_0_660 (.ZN (\partial_reg[19][0] ), .A1 (n_4_0_51), .A2 (n_4_0_1));
INV_X2 i_4_0_659 (.ZN (n_4_0_51), .A (\op2[19] ));
NOR2_X1 i_4_0_658 (.ZN (\partial_reg[18][31] ), .A1 (n_4_0_50), .A2 (n_4_0_32));
NOR2_X1 i_4_0_657 (.ZN (\partial_reg[18][30] ), .A1 (n_4_0_50), .A2 (n_4_0_31));
NOR2_X1 i_4_0_656 (.ZN (\partial_reg[18][29] ), .A1 (n_4_0_50), .A2 (n_4_0_30));
NOR2_X1 i_4_0_655 (.ZN (\partial_reg[18][28] ), .A1 (n_4_0_50), .A2 (n_4_0_29));
NOR2_X1 i_4_0_654 (.ZN (\partial_reg[18][27] ), .A1 (n_4_0_50), .A2 (n_4_0_28));
NOR2_X1 i_4_0_653 (.ZN (\partial_reg[18][26] ), .A1 (n_4_0_50), .A2 (n_4_0_27));
NOR2_X1 i_4_0_652 (.ZN (\partial_reg[18][25] ), .A1 (n_4_0_50), .A2 (n_4_0_26));
NOR2_X1 i_4_0_651 (.ZN (\partial_reg[18][24] ), .A1 (n_4_0_50), .A2 (n_4_0_25));
NOR2_X1 i_4_0_650 (.ZN (\partial_reg[18][23] ), .A1 (n_4_0_50), .A2 (n_4_0_24));
NOR2_X1 i_4_0_649 (.ZN (\partial_reg[18][22] ), .A1 (n_4_0_50), .A2 (n_4_0_23));
NOR2_X1 i_4_0_648 (.ZN (\partial_reg[18][21] ), .A1 (n_4_0_50), .A2 (n_4_0_22));
NOR2_X1 i_4_0_647 (.ZN (\partial_reg[18][20] ), .A1 (n_4_0_50), .A2 (n_4_0_21));
NOR2_X1 i_4_0_646 (.ZN (\partial_reg[18][19] ), .A1 (n_4_0_50), .A2 (n_4_0_20));
NOR2_X1 i_4_0_645 (.ZN (\partial_reg[18][18] ), .A1 (n_4_0_50), .A2 (n_4_0_19));
NOR2_X1 i_4_0_644 (.ZN (\partial_reg[18][17] ), .A1 (n_4_0_50), .A2 (n_4_0_18));
NOR2_X1 i_4_0_643 (.ZN (\partial_reg[18][16] ), .A1 (n_4_0_50), .A2 (n_4_0_17));
NOR2_X1 i_4_0_642 (.ZN (\partial_reg[18][15] ), .A1 (n_4_0_50), .A2 (n_4_0_16));
NOR2_X1 i_4_0_641 (.ZN (\partial_reg[18][14] ), .A1 (n_4_0_50), .A2 (n_4_0_15));
NOR2_X1 i_4_0_640 (.ZN (\partial_reg[18][13] ), .A1 (n_4_0_50), .A2 (n_4_0_14));
NOR2_X1 i_4_0_639 (.ZN (\partial_reg[18][12] ), .A1 (n_4_0_50), .A2 (n_4_0_13));
NOR2_X1 i_4_0_638 (.ZN (\partial_reg[18][11] ), .A1 (n_4_0_50), .A2 (n_4_0_12));
NOR2_X1 i_4_0_637 (.ZN (\partial_reg[18][10] ), .A1 (n_4_0_50), .A2 (n_4_0_11));
NOR2_X1 i_4_0_636 (.ZN (\partial_reg[18][9] ), .A1 (n_4_0_50), .A2 (n_4_0_10));
NOR2_X1 i_4_0_635 (.ZN (\partial_reg[18][8] ), .A1 (n_4_0_50), .A2 (n_4_0_9));
NOR2_X1 i_4_0_634 (.ZN (\partial_reg[18][7] ), .A1 (n_4_0_50), .A2 (n_4_0_8));
NOR2_X1 i_4_0_633 (.ZN (\partial_reg[18][6] ), .A1 (n_4_0_50), .A2 (n_4_0_7));
NOR2_X1 i_4_0_632 (.ZN (\partial_reg[18][5] ), .A1 (n_4_0_50), .A2 (n_4_0_6));
NOR2_X1 i_4_0_631 (.ZN (\partial_reg[18][4] ), .A1 (n_4_0_50), .A2 (n_4_0_5));
NOR2_X1 i_4_0_630 (.ZN (\partial_reg[18][3] ), .A1 (n_4_0_50), .A2 (n_4_0_4));
NOR2_X1 i_4_0_629 (.ZN (\partial_reg[18][2] ), .A1 (n_4_0_50), .A2 (n_4_0_3));
NOR2_X1 i_4_0_628 (.ZN (\partial_reg[18][1] ), .A1 (n_4_0_50), .A2 (n_4_0_2));
NOR2_X1 i_4_0_627 (.ZN (\partial_reg[18][0] ), .A1 (n_4_0_50), .A2 (n_4_0_1));
INV_X2 i_4_0_626 (.ZN (n_4_0_50), .A (\op2[18] ));
NOR2_X1 i_4_0_625 (.ZN (\partial_reg[17][31] ), .A1 (n_4_0_49), .A2 (n_4_0_32));
NOR2_X1 i_4_0_624 (.ZN (\partial_reg[17][30] ), .A1 (n_4_0_49), .A2 (n_4_0_31));
NOR2_X1 i_4_0_623 (.ZN (\partial_reg[17][29] ), .A1 (n_4_0_49), .A2 (n_4_0_30));
NOR2_X1 i_4_0_622 (.ZN (\partial_reg[17][28] ), .A1 (n_4_0_49), .A2 (n_4_0_29));
NOR2_X1 i_4_0_621 (.ZN (\partial_reg[17][27] ), .A1 (n_4_0_49), .A2 (n_4_0_28));
NOR2_X1 i_4_0_620 (.ZN (\partial_reg[17][26] ), .A1 (n_4_0_49), .A2 (n_4_0_27));
NOR2_X1 i_4_0_619 (.ZN (\partial_reg[17][25] ), .A1 (n_4_0_49), .A2 (n_4_0_26));
NOR2_X1 i_4_0_618 (.ZN (\partial_reg[17][24] ), .A1 (n_4_0_49), .A2 (n_4_0_25));
NOR2_X1 i_4_0_617 (.ZN (\partial_reg[17][23] ), .A1 (n_4_0_49), .A2 (n_4_0_24));
NOR2_X1 i_4_0_616 (.ZN (\partial_reg[17][22] ), .A1 (n_4_0_49), .A2 (n_4_0_23));
NOR2_X1 i_4_0_615 (.ZN (\partial_reg[17][21] ), .A1 (n_4_0_49), .A2 (n_4_0_22));
NOR2_X1 i_4_0_614 (.ZN (\partial_reg[17][20] ), .A1 (n_4_0_49), .A2 (n_4_0_21));
NOR2_X1 i_4_0_613 (.ZN (\partial_reg[17][19] ), .A1 (n_4_0_49), .A2 (n_4_0_20));
NOR2_X1 i_4_0_612 (.ZN (\partial_reg[17][18] ), .A1 (n_4_0_49), .A2 (n_4_0_19));
NOR2_X1 i_4_0_611 (.ZN (\partial_reg[17][17] ), .A1 (n_4_0_49), .A2 (n_4_0_18));
NOR2_X1 i_4_0_610 (.ZN (\partial_reg[17][16] ), .A1 (n_4_0_49), .A2 (n_4_0_17));
NOR2_X1 i_4_0_609 (.ZN (\partial_reg[17][15] ), .A1 (n_4_0_49), .A2 (n_4_0_16));
NOR2_X1 i_4_0_608 (.ZN (\partial_reg[17][14] ), .A1 (n_4_0_49), .A2 (n_4_0_15));
NOR2_X1 i_4_0_607 (.ZN (\partial_reg[17][13] ), .A1 (n_4_0_49), .A2 (n_4_0_14));
NOR2_X1 i_4_0_606 (.ZN (\partial_reg[17][12] ), .A1 (n_4_0_49), .A2 (n_4_0_13));
NOR2_X1 i_4_0_605 (.ZN (\partial_reg[17][11] ), .A1 (n_4_0_49), .A2 (n_4_0_12));
NOR2_X1 i_4_0_604 (.ZN (\partial_reg[17][10] ), .A1 (n_4_0_49), .A2 (n_4_0_11));
NOR2_X1 i_4_0_603 (.ZN (\partial_reg[17][9] ), .A1 (n_4_0_49), .A2 (n_4_0_10));
NOR2_X1 i_4_0_602 (.ZN (\partial_reg[17][8] ), .A1 (n_4_0_49), .A2 (n_4_0_9));
NOR2_X1 i_4_0_601 (.ZN (\partial_reg[17][7] ), .A1 (n_4_0_49), .A2 (n_4_0_8));
NOR2_X1 i_4_0_600 (.ZN (\partial_reg[17][6] ), .A1 (n_4_0_49), .A2 (n_4_0_7));
NOR2_X1 i_4_0_599 (.ZN (\partial_reg[17][5] ), .A1 (n_4_0_49), .A2 (n_4_0_6));
NOR2_X1 i_4_0_598 (.ZN (\partial_reg[17][4] ), .A1 (n_4_0_49), .A2 (n_4_0_5));
NOR2_X1 i_4_0_597 (.ZN (\partial_reg[17][3] ), .A1 (n_4_0_49), .A2 (n_4_0_4));
NOR2_X1 i_4_0_596 (.ZN (\partial_reg[17][2] ), .A1 (n_4_0_49), .A2 (n_4_0_3));
NOR2_X1 i_4_0_595 (.ZN (\partial_reg[17][1] ), .A1 (n_4_0_49), .A2 (n_4_0_2));
NOR2_X1 i_4_0_594 (.ZN (\partial_reg[17][0] ), .A1 (n_4_0_49), .A2 (n_4_0_1));
INV_X2 i_4_0_593 (.ZN (n_4_0_49), .A (\op2[17] ));
NOR2_X1 i_4_0_592 (.ZN (\partial_reg[16][31] ), .A1 (n_4_0_48), .A2 (n_4_0_32));
NOR2_X1 i_4_0_591 (.ZN (\partial_reg[16][30] ), .A1 (n_4_0_48), .A2 (n_4_0_31));
NOR2_X1 i_4_0_590 (.ZN (\partial_reg[16][29] ), .A1 (n_4_0_48), .A2 (n_4_0_30));
NOR2_X1 i_4_0_589 (.ZN (\partial_reg[16][28] ), .A1 (n_4_0_48), .A2 (n_4_0_29));
NOR2_X1 i_4_0_588 (.ZN (\partial_reg[16][27] ), .A1 (n_4_0_48), .A2 (n_4_0_28));
NOR2_X1 i_4_0_587 (.ZN (\partial_reg[16][26] ), .A1 (n_4_0_48), .A2 (n_4_0_27));
NOR2_X1 i_4_0_586 (.ZN (\partial_reg[16][25] ), .A1 (n_4_0_48), .A2 (n_4_0_26));
NOR2_X1 i_4_0_585 (.ZN (\partial_reg[16][24] ), .A1 (n_4_0_48), .A2 (n_4_0_25));
NOR2_X1 i_4_0_584 (.ZN (\partial_reg[16][23] ), .A1 (n_4_0_48), .A2 (n_4_0_24));
NOR2_X1 i_4_0_583 (.ZN (\partial_reg[16][22] ), .A1 (n_4_0_48), .A2 (n_4_0_23));
NOR2_X1 i_4_0_582 (.ZN (\partial_reg[16][21] ), .A1 (n_4_0_48), .A2 (n_4_0_22));
NOR2_X1 i_4_0_581 (.ZN (\partial_reg[16][20] ), .A1 (n_4_0_48), .A2 (n_4_0_21));
NOR2_X1 i_4_0_580 (.ZN (\partial_reg[16][19] ), .A1 (n_4_0_48), .A2 (n_4_0_20));
NOR2_X1 i_4_0_579 (.ZN (\partial_reg[16][18] ), .A1 (n_4_0_48), .A2 (n_4_0_19));
NOR2_X1 i_4_0_578 (.ZN (\partial_reg[16][17] ), .A1 (n_4_0_48), .A2 (n_4_0_18));
NOR2_X1 i_4_0_577 (.ZN (\partial_reg[16][16] ), .A1 (n_4_0_48), .A2 (n_4_0_17));
NOR2_X1 i_4_0_576 (.ZN (\partial_reg[16][15] ), .A1 (n_4_0_48), .A2 (n_4_0_16));
NOR2_X1 i_4_0_575 (.ZN (\partial_reg[16][14] ), .A1 (n_4_0_48), .A2 (n_4_0_15));
NOR2_X1 i_4_0_574 (.ZN (\partial_reg[16][13] ), .A1 (n_4_0_48), .A2 (n_4_0_14));
NOR2_X1 i_4_0_573 (.ZN (\partial_reg[16][12] ), .A1 (n_4_0_48), .A2 (n_4_0_13));
NOR2_X1 i_4_0_572 (.ZN (\partial_reg[16][11] ), .A1 (n_4_0_48), .A2 (n_4_0_12));
NOR2_X1 i_4_0_571 (.ZN (\partial_reg[16][10] ), .A1 (n_4_0_48), .A2 (n_4_0_11));
NOR2_X1 i_4_0_570 (.ZN (\partial_reg[16][9] ), .A1 (n_4_0_48), .A2 (n_4_0_10));
NOR2_X1 i_4_0_569 (.ZN (\partial_reg[16][8] ), .A1 (n_4_0_48), .A2 (n_4_0_9));
NOR2_X1 i_4_0_568 (.ZN (\partial_reg[16][7] ), .A1 (n_4_0_48), .A2 (n_4_0_8));
NOR2_X1 i_4_0_567 (.ZN (\partial_reg[16][6] ), .A1 (n_4_0_48), .A2 (n_4_0_7));
NOR2_X1 i_4_0_566 (.ZN (\partial_reg[16][5] ), .A1 (n_4_0_48), .A2 (n_4_0_6));
NOR2_X1 i_4_0_565 (.ZN (\partial_reg[16][4] ), .A1 (n_4_0_48), .A2 (n_4_0_5));
NOR2_X1 i_4_0_564 (.ZN (\partial_reg[16][3] ), .A1 (n_4_0_48), .A2 (n_4_0_4));
NOR2_X1 i_4_0_563 (.ZN (\partial_reg[16][2] ), .A1 (n_4_0_48), .A2 (n_4_0_3));
NOR2_X1 i_4_0_562 (.ZN (\partial_reg[16][1] ), .A1 (n_4_0_48), .A2 (n_4_0_2));
NOR2_X1 i_4_0_561 (.ZN (\partial_reg[16][0] ), .A1 (n_4_0_48), .A2 (n_4_0_1));
INV_X2 i_4_0_560 (.ZN (n_4_0_48), .A (\op2[16] ));
NOR2_X1 i_4_0_559 (.ZN (\partial_reg[15][31] ), .A1 (n_4_0_47), .A2 (n_4_0_32));
NOR2_X1 i_4_0_558 (.ZN (\partial_reg[15][30] ), .A1 (n_4_0_47), .A2 (n_4_0_31));
NOR2_X1 i_4_0_557 (.ZN (\partial_reg[15][29] ), .A1 (n_4_0_47), .A2 (n_4_0_30));
NOR2_X1 i_4_0_556 (.ZN (\partial_reg[15][28] ), .A1 (n_4_0_47), .A2 (n_4_0_29));
NOR2_X1 i_4_0_555 (.ZN (\partial_reg[15][27] ), .A1 (n_4_0_47), .A2 (n_4_0_28));
NOR2_X1 i_4_0_554 (.ZN (\partial_reg[15][26] ), .A1 (n_4_0_47), .A2 (n_4_0_27));
NOR2_X1 i_4_0_553 (.ZN (\partial_reg[15][25] ), .A1 (n_4_0_47), .A2 (n_4_0_26));
NOR2_X1 i_4_0_552 (.ZN (\partial_reg[15][24] ), .A1 (n_4_0_47), .A2 (n_4_0_25));
NOR2_X1 i_4_0_551 (.ZN (\partial_reg[15][23] ), .A1 (n_4_0_47), .A2 (n_4_0_24));
NOR2_X1 i_4_0_550 (.ZN (\partial_reg[15][22] ), .A1 (n_4_0_47), .A2 (n_4_0_23));
NOR2_X1 i_4_0_549 (.ZN (\partial_reg[15][21] ), .A1 (n_4_0_47), .A2 (n_4_0_22));
NOR2_X1 i_4_0_548 (.ZN (\partial_reg[15][20] ), .A1 (n_4_0_47), .A2 (n_4_0_21));
NOR2_X1 i_4_0_547 (.ZN (\partial_reg[15][19] ), .A1 (n_4_0_47), .A2 (n_4_0_20));
NOR2_X1 i_4_0_546 (.ZN (\partial_reg[15][18] ), .A1 (n_4_0_47), .A2 (n_4_0_19));
NOR2_X1 i_4_0_545 (.ZN (\partial_reg[15][17] ), .A1 (n_4_0_47), .A2 (n_4_0_18));
NOR2_X1 i_4_0_544 (.ZN (\partial_reg[15][16] ), .A1 (n_4_0_47), .A2 (n_4_0_17));
NOR2_X1 i_4_0_543 (.ZN (\partial_reg[15][15] ), .A1 (n_4_0_47), .A2 (n_4_0_16));
NOR2_X1 i_4_0_542 (.ZN (\partial_reg[15][14] ), .A1 (n_4_0_47), .A2 (n_4_0_15));
NOR2_X1 i_4_0_541 (.ZN (\partial_reg[15][13] ), .A1 (n_4_0_47), .A2 (n_4_0_14));
NOR2_X1 i_4_0_540 (.ZN (\partial_reg[15][12] ), .A1 (n_4_0_47), .A2 (n_4_0_13));
NOR2_X1 i_4_0_539 (.ZN (\partial_reg[15][11] ), .A1 (n_4_0_47), .A2 (n_4_0_12));
NOR2_X1 i_4_0_538 (.ZN (\partial_reg[15][10] ), .A1 (n_4_0_47), .A2 (n_4_0_11));
NOR2_X1 i_4_0_537 (.ZN (\partial_reg[15][9] ), .A1 (n_4_0_47), .A2 (n_4_0_10));
NOR2_X1 i_4_0_536 (.ZN (\partial_reg[15][8] ), .A1 (n_4_0_47), .A2 (n_4_0_9));
NOR2_X1 i_4_0_535 (.ZN (\partial_reg[15][7] ), .A1 (n_4_0_47), .A2 (n_4_0_8));
NOR2_X1 i_4_0_534 (.ZN (\partial_reg[15][6] ), .A1 (n_4_0_47), .A2 (n_4_0_7));
NOR2_X1 i_4_0_533 (.ZN (\partial_reg[15][5] ), .A1 (n_4_0_47), .A2 (n_4_0_6));
NOR2_X1 i_4_0_532 (.ZN (\partial_reg[15][4] ), .A1 (n_4_0_47), .A2 (n_4_0_5));
NOR2_X1 i_4_0_531 (.ZN (\partial_reg[15][3] ), .A1 (n_4_0_47), .A2 (n_4_0_4));
NOR2_X1 i_4_0_530 (.ZN (\partial_reg[15][2] ), .A1 (n_4_0_47), .A2 (n_4_0_3));
NOR2_X1 i_4_0_529 (.ZN (\partial_reg[15][1] ), .A1 (n_4_0_47), .A2 (n_4_0_2));
NOR2_X1 i_4_0_528 (.ZN (\partial_reg[15][0] ), .A1 (n_4_0_47), .A2 (n_4_0_1));
INV_X2 i_4_0_527 (.ZN (n_4_0_47), .A (\op2[15] ));
NOR2_X1 i_4_0_526 (.ZN (\partial_reg[14][31] ), .A1 (n_4_0_46), .A2 (n_4_0_32));
NOR2_X1 i_4_0_525 (.ZN (\partial_reg[14][30] ), .A1 (n_4_0_46), .A2 (n_4_0_31));
NOR2_X1 i_4_0_524 (.ZN (\partial_reg[14][29] ), .A1 (n_4_0_46), .A2 (n_4_0_30));
NOR2_X1 i_4_0_523 (.ZN (\partial_reg[14][28] ), .A1 (n_4_0_46), .A2 (n_4_0_29));
NOR2_X1 i_4_0_522 (.ZN (\partial_reg[14][27] ), .A1 (n_4_0_46), .A2 (n_4_0_28));
NOR2_X1 i_4_0_521 (.ZN (\partial_reg[14][26] ), .A1 (n_4_0_46), .A2 (n_4_0_27));
NOR2_X1 i_4_0_520 (.ZN (\partial_reg[14][25] ), .A1 (n_4_0_46), .A2 (n_4_0_26));
NOR2_X1 i_4_0_519 (.ZN (\partial_reg[14][24] ), .A1 (n_4_0_46), .A2 (n_4_0_25));
NOR2_X1 i_4_0_518 (.ZN (\partial_reg[14][23] ), .A1 (n_4_0_46), .A2 (n_4_0_24));
NOR2_X1 i_4_0_517 (.ZN (\partial_reg[14][22] ), .A1 (n_4_0_46), .A2 (n_4_0_23));
NOR2_X1 i_4_0_516 (.ZN (\partial_reg[14][21] ), .A1 (n_4_0_46), .A2 (n_4_0_22));
NOR2_X1 i_4_0_515 (.ZN (\partial_reg[14][20] ), .A1 (n_4_0_46), .A2 (n_4_0_21));
NOR2_X1 i_4_0_514 (.ZN (\partial_reg[14][19] ), .A1 (n_4_0_46), .A2 (n_4_0_20));
NOR2_X1 i_4_0_513 (.ZN (\partial_reg[14][18] ), .A1 (n_4_0_46), .A2 (n_4_0_19));
NOR2_X1 i_4_0_512 (.ZN (\partial_reg[14][17] ), .A1 (n_4_0_46), .A2 (n_4_0_18));
NOR2_X1 i_4_0_511 (.ZN (\partial_reg[14][16] ), .A1 (n_4_0_46), .A2 (n_4_0_17));
NOR2_X1 i_4_0_510 (.ZN (\partial_reg[14][15] ), .A1 (n_4_0_46), .A2 (n_4_0_16));
NOR2_X1 i_4_0_509 (.ZN (\partial_reg[14][14] ), .A1 (n_4_0_46), .A2 (n_4_0_15));
NOR2_X1 i_4_0_508 (.ZN (\partial_reg[14][13] ), .A1 (n_4_0_46), .A2 (n_4_0_14));
NOR2_X1 i_4_0_507 (.ZN (\partial_reg[14][12] ), .A1 (n_4_0_46), .A2 (n_4_0_13));
NOR2_X1 i_4_0_506 (.ZN (\partial_reg[14][11] ), .A1 (n_4_0_46), .A2 (n_4_0_12));
NOR2_X1 i_4_0_505 (.ZN (\partial_reg[14][10] ), .A1 (n_4_0_46), .A2 (n_4_0_11));
NOR2_X1 i_4_0_504 (.ZN (\partial_reg[14][9] ), .A1 (n_4_0_46), .A2 (n_4_0_10));
NOR2_X1 i_4_0_503 (.ZN (\partial_reg[14][8] ), .A1 (n_4_0_46), .A2 (n_4_0_9));
NOR2_X1 i_4_0_502 (.ZN (\partial_reg[14][7] ), .A1 (n_4_0_46), .A2 (n_4_0_8));
NOR2_X1 i_4_0_501 (.ZN (\partial_reg[14][6] ), .A1 (n_4_0_46), .A2 (n_4_0_7));
NOR2_X1 i_4_0_500 (.ZN (\partial_reg[14][5] ), .A1 (n_4_0_46), .A2 (n_4_0_6));
NOR2_X1 i_4_0_499 (.ZN (\partial_reg[14][4] ), .A1 (n_4_0_46), .A2 (n_4_0_5));
NOR2_X1 i_4_0_498 (.ZN (\partial_reg[14][3] ), .A1 (n_4_0_46), .A2 (n_4_0_4));
NOR2_X1 i_4_0_497 (.ZN (\partial_reg[14][2] ), .A1 (n_4_0_46), .A2 (n_4_0_3));
NOR2_X1 i_4_0_496 (.ZN (\partial_reg[14][1] ), .A1 (n_4_0_46), .A2 (n_4_0_2));
NOR2_X1 i_4_0_495 (.ZN (\partial_reg[14][0] ), .A1 (n_4_0_46), .A2 (n_4_0_1));
INV_X2 i_4_0_494 (.ZN (n_4_0_46), .A (\op2[14] ));
NOR2_X1 i_4_0_493 (.ZN (\partial_reg[13][31] ), .A1 (n_4_0_45), .A2 (n_4_0_32));
NOR2_X1 i_4_0_492 (.ZN (\partial_reg[13][30] ), .A1 (n_4_0_45), .A2 (n_4_0_31));
NOR2_X1 i_4_0_491 (.ZN (\partial_reg[13][29] ), .A1 (n_4_0_45), .A2 (n_4_0_30));
NOR2_X1 i_4_0_490 (.ZN (\partial_reg[13][28] ), .A1 (n_4_0_45), .A2 (n_4_0_29));
NOR2_X1 i_4_0_489 (.ZN (\partial_reg[13][27] ), .A1 (n_4_0_45), .A2 (n_4_0_28));
NOR2_X1 i_4_0_488 (.ZN (\partial_reg[13][26] ), .A1 (n_4_0_45), .A2 (n_4_0_27));
NOR2_X1 i_4_0_487 (.ZN (\partial_reg[13][25] ), .A1 (n_4_0_45), .A2 (n_4_0_26));
NOR2_X1 i_4_0_486 (.ZN (\partial_reg[13][24] ), .A1 (n_4_0_45), .A2 (n_4_0_25));
NOR2_X1 i_4_0_485 (.ZN (\partial_reg[13][23] ), .A1 (n_4_0_45), .A2 (n_4_0_24));
NOR2_X1 i_4_0_484 (.ZN (\partial_reg[13][22] ), .A1 (n_4_0_45), .A2 (n_4_0_23));
NOR2_X1 i_4_0_483 (.ZN (\partial_reg[13][21] ), .A1 (n_4_0_45), .A2 (n_4_0_22));
NOR2_X1 i_4_0_482 (.ZN (\partial_reg[13][20] ), .A1 (n_4_0_45), .A2 (n_4_0_21));
NOR2_X1 i_4_0_481 (.ZN (\partial_reg[13][19] ), .A1 (n_4_0_45), .A2 (n_4_0_20));
NOR2_X1 i_4_0_480 (.ZN (\partial_reg[13][18] ), .A1 (n_4_0_45), .A2 (n_4_0_19));
NOR2_X1 i_4_0_479 (.ZN (\partial_reg[13][17] ), .A1 (n_4_0_45), .A2 (n_4_0_18));
NOR2_X1 i_4_0_478 (.ZN (\partial_reg[13][16] ), .A1 (n_4_0_45), .A2 (n_4_0_17));
NOR2_X1 i_4_0_477 (.ZN (\partial_reg[13][15] ), .A1 (n_4_0_45), .A2 (n_4_0_16));
NOR2_X1 i_4_0_476 (.ZN (\partial_reg[13][14] ), .A1 (n_4_0_45), .A2 (n_4_0_15));
NOR2_X1 i_4_0_475 (.ZN (\partial_reg[13][13] ), .A1 (n_4_0_45), .A2 (n_4_0_14));
NOR2_X1 i_4_0_474 (.ZN (\partial_reg[13][12] ), .A1 (n_4_0_45), .A2 (n_4_0_13));
NOR2_X1 i_4_0_473 (.ZN (\partial_reg[13][11] ), .A1 (n_4_0_45), .A2 (n_4_0_12));
NOR2_X1 i_4_0_472 (.ZN (\partial_reg[13][10] ), .A1 (n_4_0_45), .A2 (n_4_0_11));
NOR2_X1 i_4_0_471 (.ZN (\partial_reg[13][9] ), .A1 (n_4_0_45), .A2 (n_4_0_10));
NOR2_X1 i_4_0_470 (.ZN (\partial_reg[13][8] ), .A1 (n_4_0_45), .A2 (n_4_0_9));
NOR2_X1 i_4_0_469 (.ZN (\partial_reg[13][7] ), .A1 (n_4_0_45), .A2 (n_4_0_8));
NOR2_X1 i_4_0_468 (.ZN (\partial_reg[13][6] ), .A1 (n_4_0_45), .A2 (n_4_0_7));
NOR2_X1 i_4_0_467 (.ZN (\partial_reg[13][5] ), .A1 (n_4_0_45), .A2 (n_4_0_6));
NOR2_X1 i_4_0_466 (.ZN (\partial_reg[13][4] ), .A1 (n_4_0_45), .A2 (n_4_0_5));
NOR2_X1 i_4_0_465 (.ZN (\partial_reg[13][3] ), .A1 (n_4_0_45), .A2 (n_4_0_4));
NOR2_X1 i_4_0_464 (.ZN (\partial_reg[13][2] ), .A1 (n_4_0_45), .A2 (n_4_0_3));
NOR2_X1 i_4_0_463 (.ZN (\partial_reg[13][1] ), .A1 (n_4_0_45), .A2 (n_4_0_2));
NOR2_X1 i_4_0_462 (.ZN (\partial_reg[13][0] ), .A1 (n_4_0_45), .A2 (n_4_0_1));
INV_X2 i_4_0_461 (.ZN (n_4_0_45), .A (\op2[13] ));
NOR2_X1 i_4_0_460 (.ZN (\partial_reg[12][31] ), .A1 (n_4_0_44), .A2 (n_4_0_32));
NOR2_X1 i_4_0_459 (.ZN (\partial_reg[12][30] ), .A1 (n_4_0_44), .A2 (n_4_0_31));
NOR2_X1 i_4_0_458 (.ZN (\partial_reg[12][29] ), .A1 (n_4_0_44), .A2 (n_4_0_30));
NOR2_X1 i_4_0_457 (.ZN (\partial_reg[12][28] ), .A1 (n_4_0_44), .A2 (n_4_0_29));
NOR2_X1 i_4_0_456 (.ZN (\partial_reg[12][27] ), .A1 (n_4_0_44), .A2 (n_4_0_28));
NOR2_X1 i_4_0_455 (.ZN (\partial_reg[12][26] ), .A1 (n_4_0_44), .A2 (n_4_0_27));
NOR2_X1 i_4_0_454 (.ZN (\partial_reg[12][25] ), .A1 (n_4_0_44), .A2 (n_4_0_26));
NOR2_X1 i_4_0_453 (.ZN (\partial_reg[12][24] ), .A1 (n_4_0_44), .A2 (n_4_0_25));
NOR2_X1 i_4_0_452 (.ZN (\partial_reg[12][23] ), .A1 (n_4_0_44), .A2 (n_4_0_24));
NOR2_X1 i_4_0_451 (.ZN (\partial_reg[12][22] ), .A1 (n_4_0_44), .A2 (n_4_0_23));
NOR2_X1 i_4_0_450 (.ZN (\partial_reg[12][21] ), .A1 (n_4_0_44), .A2 (n_4_0_22));
NOR2_X1 i_4_0_449 (.ZN (\partial_reg[12][20] ), .A1 (n_4_0_44), .A2 (n_4_0_21));
NOR2_X1 i_4_0_448 (.ZN (\partial_reg[12][19] ), .A1 (n_4_0_44), .A2 (n_4_0_20));
NOR2_X1 i_4_0_447 (.ZN (\partial_reg[12][18] ), .A1 (n_4_0_44), .A2 (n_4_0_19));
NOR2_X1 i_4_0_446 (.ZN (\partial_reg[12][17] ), .A1 (n_4_0_44), .A2 (n_4_0_18));
NOR2_X1 i_4_0_445 (.ZN (\partial_reg[12][16] ), .A1 (n_4_0_44), .A2 (n_4_0_17));
NOR2_X1 i_4_0_444 (.ZN (\partial_reg[12][15] ), .A1 (n_4_0_44), .A2 (n_4_0_16));
NOR2_X1 i_4_0_443 (.ZN (\partial_reg[12][14] ), .A1 (n_4_0_44), .A2 (n_4_0_15));
NOR2_X1 i_4_0_442 (.ZN (\partial_reg[12][13] ), .A1 (n_4_0_44), .A2 (n_4_0_14));
NOR2_X1 i_4_0_441 (.ZN (\partial_reg[12][12] ), .A1 (n_4_0_44), .A2 (n_4_0_13));
NOR2_X1 i_4_0_440 (.ZN (\partial_reg[12][11] ), .A1 (n_4_0_44), .A2 (n_4_0_12));
NOR2_X1 i_4_0_439 (.ZN (\partial_reg[12][10] ), .A1 (n_4_0_44), .A2 (n_4_0_11));
NOR2_X1 i_4_0_438 (.ZN (\partial_reg[12][9] ), .A1 (n_4_0_44), .A2 (n_4_0_10));
NOR2_X1 i_4_0_437 (.ZN (\partial_reg[12][8] ), .A1 (n_4_0_44), .A2 (n_4_0_9));
NOR2_X1 i_4_0_436 (.ZN (\partial_reg[12][7] ), .A1 (n_4_0_44), .A2 (n_4_0_8));
NOR2_X1 i_4_0_435 (.ZN (\partial_reg[12][6] ), .A1 (n_4_0_44), .A2 (n_4_0_7));
NOR2_X1 i_4_0_434 (.ZN (\partial_reg[12][5] ), .A1 (n_4_0_44), .A2 (n_4_0_6));
NOR2_X1 i_4_0_433 (.ZN (\partial_reg[12][4] ), .A1 (n_4_0_44), .A2 (n_4_0_5));
NOR2_X1 i_4_0_432 (.ZN (\partial_reg[12][3] ), .A1 (n_4_0_44), .A2 (n_4_0_4));
NOR2_X1 i_4_0_431 (.ZN (\partial_reg[12][2] ), .A1 (n_4_0_44), .A2 (n_4_0_3));
NOR2_X1 i_4_0_430 (.ZN (\partial_reg[12][1] ), .A1 (n_4_0_44), .A2 (n_4_0_2));
NOR2_X1 i_4_0_429 (.ZN (\partial_reg[12][0] ), .A1 (n_4_0_44), .A2 (n_4_0_1));
INV_X2 i_4_0_428 (.ZN (n_4_0_44), .A (\op2[12] ));
NOR2_X1 i_4_0_427 (.ZN (\partial_reg[11][31] ), .A1 (n_4_0_43), .A2 (n_4_0_32));
NOR2_X1 i_4_0_426 (.ZN (\partial_reg[11][30] ), .A1 (n_4_0_43), .A2 (n_4_0_31));
NOR2_X1 i_4_0_425 (.ZN (\partial_reg[11][29] ), .A1 (n_4_0_43), .A2 (n_4_0_30));
NOR2_X1 i_4_0_424 (.ZN (\partial_reg[11][28] ), .A1 (n_4_0_43), .A2 (n_4_0_29));
NOR2_X1 i_4_0_423 (.ZN (\partial_reg[11][27] ), .A1 (n_4_0_43), .A2 (n_4_0_28));
NOR2_X1 i_4_0_422 (.ZN (\partial_reg[11][26] ), .A1 (n_4_0_43), .A2 (n_4_0_27));
NOR2_X1 i_4_0_421 (.ZN (\partial_reg[11][25] ), .A1 (n_4_0_43), .A2 (n_4_0_26));
NOR2_X1 i_4_0_420 (.ZN (\partial_reg[11][24] ), .A1 (n_4_0_43), .A2 (n_4_0_25));
NOR2_X1 i_4_0_419 (.ZN (\partial_reg[11][23] ), .A1 (n_4_0_43), .A2 (n_4_0_24));
NOR2_X1 i_4_0_418 (.ZN (\partial_reg[11][22] ), .A1 (n_4_0_43), .A2 (n_4_0_23));
NOR2_X1 i_4_0_417 (.ZN (\partial_reg[11][21] ), .A1 (n_4_0_43), .A2 (n_4_0_22));
NOR2_X1 i_4_0_416 (.ZN (\partial_reg[11][20] ), .A1 (n_4_0_43), .A2 (n_4_0_21));
NOR2_X1 i_4_0_415 (.ZN (\partial_reg[11][19] ), .A1 (n_4_0_43), .A2 (n_4_0_20));
NOR2_X1 i_4_0_414 (.ZN (\partial_reg[11][18] ), .A1 (n_4_0_43), .A2 (n_4_0_19));
NOR2_X1 i_4_0_413 (.ZN (\partial_reg[11][17] ), .A1 (n_4_0_43), .A2 (n_4_0_18));
NOR2_X1 i_4_0_412 (.ZN (\partial_reg[11][16] ), .A1 (n_4_0_43), .A2 (n_4_0_17));
NOR2_X1 i_4_0_411 (.ZN (\partial_reg[11][15] ), .A1 (n_4_0_43), .A2 (n_4_0_16));
NOR2_X1 i_4_0_410 (.ZN (\partial_reg[11][14] ), .A1 (n_4_0_43), .A2 (n_4_0_15));
NOR2_X1 i_4_0_409 (.ZN (\partial_reg[11][13] ), .A1 (n_4_0_43), .A2 (n_4_0_14));
NOR2_X1 i_4_0_408 (.ZN (\partial_reg[11][12] ), .A1 (n_4_0_43), .A2 (n_4_0_13));
NOR2_X1 i_4_0_407 (.ZN (\partial_reg[11][11] ), .A1 (n_4_0_43), .A2 (n_4_0_12));
NOR2_X1 i_4_0_406 (.ZN (\partial_reg[11][10] ), .A1 (n_4_0_43), .A2 (n_4_0_11));
NOR2_X1 i_4_0_405 (.ZN (\partial_reg[11][9] ), .A1 (n_4_0_43), .A2 (n_4_0_10));
NOR2_X1 i_4_0_404 (.ZN (\partial_reg[11][8] ), .A1 (n_4_0_43), .A2 (n_4_0_9));
NOR2_X1 i_4_0_403 (.ZN (\partial_reg[11][7] ), .A1 (n_4_0_43), .A2 (n_4_0_8));
NOR2_X1 i_4_0_402 (.ZN (\partial_reg[11][6] ), .A1 (n_4_0_43), .A2 (n_4_0_7));
NOR2_X1 i_4_0_401 (.ZN (\partial_reg[11][5] ), .A1 (n_4_0_43), .A2 (n_4_0_6));
NOR2_X1 i_4_0_400 (.ZN (\partial_reg[11][4] ), .A1 (n_4_0_43), .A2 (n_4_0_5));
NOR2_X1 i_4_0_399 (.ZN (\partial_reg[11][3] ), .A1 (n_4_0_43), .A2 (n_4_0_4));
NOR2_X1 i_4_0_398 (.ZN (\partial_reg[11][2] ), .A1 (n_4_0_43), .A2 (n_4_0_3));
NOR2_X1 i_4_0_397 (.ZN (\partial_reg[11][1] ), .A1 (n_4_0_43), .A2 (n_4_0_2));
NOR2_X1 i_4_0_396 (.ZN (\partial_reg[11][0] ), .A1 (n_4_0_43), .A2 (n_4_0_1));
INV_X2 i_4_0_395 (.ZN (n_4_0_43), .A (\op2[11] ));
NOR2_X1 i_4_0_394 (.ZN (\partial_reg[10][31] ), .A1 (n_4_0_42), .A2 (n_4_0_32));
NOR2_X1 i_4_0_393 (.ZN (\partial_reg[10][30] ), .A1 (n_4_0_42), .A2 (n_4_0_31));
NOR2_X1 i_4_0_392 (.ZN (\partial_reg[10][29] ), .A1 (n_4_0_42), .A2 (n_4_0_30));
NOR2_X1 i_4_0_391 (.ZN (\partial_reg[10][28] ), .A1 (n_4_0_42), .A2 (n_4_0_29));
NOR2_X1 i_4_0_390 (.ZN (\partial_reg[10][27] ), .A1 (n_4_0_42), .A2 (n_4_0_28));
NOR2_X1 i_4_0_389 (.ZN (\partial_reg[10][26] ), .A1 (n_4_0_42), .A2 (n_4_0_27));
NOR2_X1 i_4_0_388 (.ZN (\partial_reg[10][25] ), .A1 (n_4_0_42), .A2 (n_4_0_26));
NOR2_X1 i_4_0_387 (.ZN (\partial_reg[10][24] ), .A1 (n_4_0_42), .A2 (n_4_0_25));
NOR2_X1 i_4_0_386 (.ZN (\partial_reg[10][23] ), .A1 (n_4_0_42), .A2 (n_4_0_24));
NOR2_X1 i_4_0_385 (.ZN (\partial_reg[10][22] ), .A1 (n_4_0_42), .A2 (n_4_0_23));
NOR2_X1 i_4_0_384 (.ZN (\partial_reg[10][21] ), .A1 (n_4_0_42), .A2 (n_4_0_22));
NOR2_X1 i_4_0_383 (.ZN (\partial_reg[10][20] ), .A1 (n_4_0_42), .A2 (n_4_0_21));
NOR2_X1 i_4_0_382 (.ZN (\partial_reg[10][19] ), .A1 (n_4_0_42), .A2 (n_4_0_20));
NOR2_X1 i_4_0_381 (.ZN (\partial_reg[10][18] ), .A1 (n_4_0_42), .A2 (n_4_0_19));
NOR2_X1 i_4_0_380 (.ZN (\partial_reg[10][17] ), .A1 (n_4_0_42), .A2 (n_4_0_18));
NOR2_X1 i_4_0_379 (.ZN (\partial_reg[10][16] ), .A1 (n_4_0_42), .A2 (n_4_0_17));
NOR2_X1 i_4_0_378 (.ZN (\partial_reg[10][15] ), .A1 (n_4_0_42), .A2 (n_4_0_16));
NOR2_X1 i_4_0_377 (.ZN (\partial_reg[10][14] ), .A1 (n_4_0_42), .A2 (n_4_0_15));
NOR2_X1 i_4_0_376 (.ZN (\partial_reg[10][13] ), .A1 (n_4_0_42), .A2 (n_4_0_14));
NOR2_X1 i_4_0_375 (.ZN (\partial_reg[10][12] ), .A1 (n_4_0_42), .A2 (n_4_0_13));
NOR2_X1 i_4_0_374 (.ZN (\partial_reg[10][11] ), .A1 (n_4_0_42), .A2 (n_4_0_12));
NOR2_X1 i_4_0_373 (.ZN (\partial_reg[10][10] ), .A1 (n_4_0_42), .A2 (n_4_0_11));
NOR2_X1 i_4_0_372 (.ZN (\partial_reg[10][9] ), .A1 (n_4_0_42), .A2 (n_4_0_10));
NOR2_X1 i_4_0_371 (.ZN (\partial_reg[10][8] ), .A1 (n_4_0_42), .A2 (n_4_0_9));
NOR2_X1 i_4_0_370 (.ZN (\partial_reg[10][7] ), .A1 (n_4_0_42), .A2 (n_4_0_8));
NOR2_X1 i_4_0_369 (.ZN (\partial_reg[10][6] ), .A1 (n_4_0_42), .A2 (n_4_0_7));
NOR2_X1 i_4_0_368 (.ZN (\partial_reg[10][5] ), .A1 (n_4_0_42), .A2 (n_4_0_6));
NOR2_X1 i_4_0_367 (.ZN (\partial_reg[10][4] ), .A1 (n_4_0_42), .A2 (n_4_0_5));
NOR2_X1 i_4_0_366 (.ZN (\partial_reg[10][3] ), .A1 (n_4_0_42), .A2 (n_4_0_4));
NOR2_X1 i_4_0_365 (.ZN (\partial_reg[10][2] ), .A1 (n_4_0_42), .A2 (n_4_0_3));
NOR2_X1 i_4_0_364 (.ZN (\partial_reg[10][1] ), .A1 (n_4_0_42), .A2 (n_4_0_2));
NOR2_X1 i_4_0_363 (.ZN (\partial_reg[10][0] ), .A1 (n_4_0_42), .A2 (n_4_0_1));
INV_X2 i_4_0_362 (.ZN (n_4_0_42), .A (\op2[10] ));
NOR2_X1 i_4_0_361 (.ZN (\partial_reg[9][31] ), .A1 (n_4_0_41), .A2 (n_4_0_32));
NOR2_X1 i_4_0_360 (.ZN (\partial_reg[9][30] ), .A1 (n_4_0_41), .A2 (n_4_0_31));
NOR2_X1 i_4_0_359 (.ZN (\partial_reg[9][29] ), .A1 (n_4_0_41), .A2 (n_4_0_30));
NOR2_X1 i_4_0_358 (.ZN (\partial_reg[9][28] ), .A1 (n_4_0_41), .A2 (n_4_0_29));
NOR2_X1 i_4_0_357 (.ZN (\partial_reg[9][27] ), .A1 (n_4_0_41), .A2 (n_4_0_28));
NOR2_X1 i_4_0_356 (.ZN (\partial_reg[9][26] ), .A1 (n_4_0_41), .A2 (n_4_0_27));
NOR2_X1 i_4_0_355 (.ZN (\partial_reg[9][25] ), .A1 (n_4_0_41), .A2 (n_4_0_26));
NOR2_X1 i_4_0_354 (.ZN (\partial_reg[9][24] ), .A1 (n_4_0_41), .A2 (n_4_0_25));
NOR2_X1 i_4_0_353 (.ZN (\partial_reg[9][23] ), .A1 (n_4_0_41), .A2 (n_4_0_24));
NOR2_X1 i_4_0_352 (.ZN (\partial_reg[9][22] ), .A1 (n_4_0_41), .A2 (n_4_0_23));
NOR2_X1 i_4_0_351 (.ZN (\partial_reg[9][21] ), .A1 (n_4_0_41), .A2 (n_4_0_22));
NOR2_X1 i_4_0_350 (.ZN (\partial_reg[9][20] ), .A1 (n_4_0_41), .A2 (n_4_0_21));
NOR2_X1 i_4_0_349 (.ZN (\partial_reg[9][19] ), .A1 (n_4_0_41), .A2 (n_4_0_20));
NOR2_X1 i_4_0_348 (.ZN (\partial_reg[9][18] ), .A1 (n_4_0_41), .A2 (n_4_0_19));
NOR2_X1 i_4_0_347 (.ZN (\partial_reg[9][17] ), .A1 (n_4_0_41), .A2 (n_4_0_18));
NOR2_X1 i_4_0_346 (.ZN (\partial_reg[9][16] ), .A1 (n_4_0_41), .A2 (n_4_0_17));
NOR2_X1 i_4_0_345 (.ZN (\partial_reg[9][15] ), .A1 (n_4_0_41), .A2 (n_4_0_16));
NOR2_X1 i_4_0_344 (.ZN (\partial_reg[9][14] ), .A1 (n_4_0_41), .A2 (n_4_0_15));
NOR2_X1 i_4_0_343 (.ZN (\partial_reg[9][13] ), .A1 (n_4_0_41), .A2 (n_4_0_14));
NOR2_X1 i_4_0_342 (.ZN (\partial_reg[9][12] ), .A1 (n_4_0_41), .A2 (n_4_0_13));
NOR2_X1 i_4_0_341 (.ZN (\partial_reg[9][11] ), .A1 (n_4_0_41), .A2 (n_4_0_12));
NOR2_X1 i_4_0_340 (.ZN (\partial_reg[9][10] ), .A1 (n_4_0_41), .A2 (n_4_0_11));
NOR2_X1 i_4_0_339 (.ZN (\partial_reg[9][9] ), .A1 (n_4_0_41), .A2 (n_4_0_10));
NOR2_X1 i_4_0_338 (.ZN (\partial_reg[9][8] ), .A1 (n_4_0_41), .A2 (n_4_0_9));
NOR2_X1 i_4_0_337 (.ZN (\partial_reg[9][7] ), .A1 (n_4_0_41), .A2 (n_4_0_8));
NOR2_X1 i_4_0_336 (.ZN (\partial_reg[9][6] ), .A1 (n_4_0_41), .A2 (n_4_0_7));
NOR2_X1 i_4_0_335 (.ZN (\partial_reg[9][5] ), .A1 (n_4_0_41), .A2 (n_4_0_6));
NOR2_X1 i_4_0_334 (.ZN (\partial_reg[9][4] ), .A1 (n_4_0_41), .A2 (n_4_0_5));
NOR2_X1 i_4_0_333 (.ZN (\partial_reg[9][3] ), .A1 (n_4_0_41), .A2 (n_4_0_4));
NOR2_X1 i_4_0_332 (.ZN (\partial_reg[9][2] ), .A1 (n_4_0_41), .A2 (n_4_0_3));
NOR2_X1 i_4_0_331 (.ZN (\partial_reg[9][1] ), .A1 (n_4_0_41), .A2 (n_4_0_2));
NOR2_X1 i_4_0_330 (.ZN (\partial_reg[9][0] ), .A1 (n_4_0_41), .A2 (n_4_0_1));
INV_X4 i_4_0_329 (.ZN (n_4_0_41), .A (\op2[9] ));
NOR2_X1 i_4_0_328 (.ZN (\partial_reg[8][31] ), .A1 (n_4_0_40), .A2 (n_4_0_32));
NOR2_X1 i_4_0_327 (.ZN (\partial_reg[8][30] ), .A1 (n_4_0_40), .A2 (n_4_0_31));
NOR2_X1 i_4_0_326 (.ZN (\partial_reg[8][29] ), .A1 (n_4_0_40), .A2 (n_4_0_30));
NOR2_X1 i_4_0_325 (.ZN (\partial_reg[8][28] ), .A1 (n_4_0_40), .A2 (n_4_0_29));
NOR2_X1 i_4_0_324 (.ZN (\partial_reg[8][27] ), .A1 (n_4_0_40), .A2 (n_4_0_28));
NOR2_X1 i_4_0_323 (.ZN (\partial_reg[8][26] ), .A1 (n_4_0_40), .A2 (n_4_0_27));
NOR2_X1 i_4_0_322 (.ZN (\partial_reg[8][25] ), .A1 (n_4_0_40), .A2 (n_4_0_26));
NOR2_X1 i_4_0_321 (.ZN (\partial_reg[8][24] ), .A1 (n_4_0_40), .A2 (n_4_0_25));
NOR2_X1 i_4_0_320 (.ZN (\partial_reg[8][23] ), .A1 (n_4_0_40), .A2 (n_4_0_24));
NOR2_X1 i_4_0_319 (.ZN (\partial_reg[8][22] ), .A1 (n_4_0_40), .A2 (n_4_0_23));
NOR2_X1 i_4_0_318 (.ZN (\partial_reg[8][21] ), .A1 (n_4_0_40), .A2 (n_4_0_22));
NOR2_X1 i_4_0_317 (.ZN (\partial_reg[8][20] ), .A1 (n_4_0_40), .A2 (n_4_0_21));
NOR2_X1 i_4_0_316 (.ZN (\partial_reg[8][19] ), .A1 (n_4_0_40), .A2 (n_4_0_20));
NOR2_X1 i_4_0_315 (.ZN (\partial_reg[8][18] ), .A1 (n_4_0_40), .A2 (n_4_0_19));
NOR2_X1 i_4_0_314 (.ZN (\partial_reg[8][17] ), .A1 (n_4_0_40), .A2 (n_4_0_18));
NOR2_X2 i_4_0_313 (.ZN (\partial_reg[8][16] ), .A1 (n_4_0_40), .A2 (n_4_0_17));
NOR2_X1 i_4_0_312 (.ZN (\partial_reg[8][15] ), .A1 (n_4_0_40), .A2 (n_4_0_16));
NOR2_X1 i_4_0_311 (.ZN (\partial_reg[8][14] ), .A1 (n_4_0_40), .A2 (n_4_0_15));
NOR2_X1 i_4_0_310 (.ZN (\partial_reg[8][13] ), .A1 (n_4_0_40), .A2 (n_4_0_14));
NOR2_X1 i_4_0_309 (.ZN (\partial_reg[8][12] ), .A1 (n_4_0_40), .A2 (n_4_0_13));
NOR2_X1 i_4_0_308 (.ZN (\partial_reg[8][11] ), .A1 (n_4_0_40), .A2 (n_4_0_12));
NOR2_X1 i_4_0_307 (.ZN (\partial_reg[8][10] ), .A1 (n_4_0_40), .A2 (n_4_0_11));
NOR2_X1 i_4_0_306 (.ZN (\partial_reg[8][9] ), .A1 (n_4_0_40), .A2 (n_4_0_10));
NOR2_X1 i_4_0_305 (.ZN (\partial_reg[8][8] ), .A1 (n_4_0_40), .A2 (n_4_0_9));
NOR2_X1 i_4_0_304 (.ZN (\partial_reg[8][7] ), .A1 (n_4_0_40), .A2 (n_4_0_8));
NOR2_X1 i_4_0_303 (.ZN (\partial_reg[8][6] ), .A1 (n_4_0_40), .A2 (n_4_0_7));
NOR2_X1 i_4_0_302 (.ZN (\partial_reg[8][5] ), .A1 (n_4_0_40), .A2 (n_4_0_6));
NOR2_X1 i_4_0_301 (.ZN (\partial_reg[8][4] ), .A1 (n_4_0_40), .A2 (n_4_0_5));
NOR2_X1 i_4_0_300 (.ZN (\partial_reg[8][3] ), .A1 (n_4_0_40), .A2 (n_4_0_4));
NOR2_X1 i_4_0_299 (.ZN (\partial_reg[8][2] ), .A1 (n_4_0_40), .A2 (n_4_0_3));
NOR2_X1 i_4_0_298 (.ZN (\partial_reg[8][1] ), .A1 (n_4_0_40), .A2 (n_4_0_2));
NOR2_X1 i_4_0_297 (.ZN (\partial_reg[8][0] ), .A1 (n_4_0_40), .A2 (n_4_0_1));
INV_X4 i_4_0_296 (.ZN (n_4_0_40), .A (\op2[8] ));
NOR2_X1 i_4_0_295 (.ZN (\partial_reg[7][31] ), .A1 (n_4_0_39), .A2 (n_4_0_32));
NOR2_X1 i_4_0_294 (.ZN (\partial_reg[7][30] ), .A1 (n_4_0_39), .A2 (n_4_0_31));
NOR2_X1 i_4_0_293 (.ZN (\partial_reg[7][29] ), .A1 (n_4_0_39), .A2 (n_4_0_30));
NOR2_X1 i_4_0_292 (.ZN (\partial_reg[7][28] ), .A1 (n_4_0_39), .A2 (n_4_0_29));
NOR2_X1 i_4_0_291 (.ZN (\partial_reg[7][27] ), .A1 (n_4_0_39), .A2 (n_4_0_28));
NOR2_X1 i_4_0_290 (.ZN (\partial_reg[7][26] ), .A1 (n_4_0_39), .A2 (n_4_0_27));
NOR2_X1 i_4_0_289 (.ZN (\partial_reg[7][25] ), .A1 (n_4_0_39), .A2 (n_4_0_26));
NOR2_X1 i_4_0_288 (.ZN (\partial_reg[7][24] ), .A1 (n_4_0_39), .A2 (n_4_0_25));
NOR2_X1 i_4_0_287 (.ZN (\partial_reg[7][23] ), .A1 (n_4_0_39), .A2 (n_4_0_24));
NOR2_X1 i_4_0_286 (.ZN (\partial_reg[7][22] ), .A1 (n_4_0_39), .A2 (n_4_0_23));
NOR2_X1 i_4_0_285 (.ZN (\partial_reg[7][21] ), .A1 (n_4_0_39), .A2 (n_4_0_22));
NOR2_X1 i_4_0_284 (.ZN (\partial_reg[7][20] ), .A1 (n_4_0_39), .A2 (n_4_0_21));
NOR2_X1 i_4_0_283 (.ZN (\partial_reg[7][19] ), .A1 (n_4_0_39), .A2 (n_4_0_20));
NOR2_X1 i_4_0_282 (.ZN (\partial_reg[7][18] ), .A1 (n_4_0_39), .A2 (n_4_0_19));
NOR2_X1 i_4_0_281 (.ZN (\partial_reg[7][17] ), .A1 (n_4_0_39), .A2 (n_4_0_18));
NOR2_X1 i_4_0_280 (.ZN (\partial_reg[7][16] ), .A1 (n_4_0_39), .A2 (n_4_0_17));
NOR2_X1 i_4_0_279 (.ZN (\partial_reg[7][15] ), .A1 (n_4_0_39), .A2 (n_4_0_16));
NOR2_X1 i_4_0_278 (.ZN (\partial_reg[7][14] ), .A1 (n_4_0_39), .A2 (n_4_0_15));
NOR2_X1 i_4_0_277 (.ZN (\partial_reg[7][13] ), .A1 (n_4_0_39), .A2 (n_4_0_14));
NOR2_X1 i_4_0_276 (.ZN (\partial_reg[7][12] ), .A1 (n_4_0_39), .A2 (n_4_0_13));
NOR2_X1 i_4_0_275 (.ZN (\partial_reg[7][11] ), .A1 (n_4_0_39), .A2 (n_4_0_12));
NOR2_X1 i_4_0_274 (.ZN (\partial_reg[7][10] ), .A1 (n_4_0_39), .A2 (n_4_0_11));
NOR2_X1 i_4_0_273 (.ZN (\partial_reg[7][9] ), .A1 (n_4_0_39), .A2 (n_4_0_10));
NOR2_X1 i_4_0_272 (.ZN (\partial_reg[7][8] ), .A1 (n_4_0_39), .A2 (n_4_0_9));
NOR2_X1 i_4_0_271 (.ZN (\partial_reg[7][7] ), .A1 (n_4_0_39), .A2 (n_4_0_8));
NOR2_X1 i_4_0_270 (.ZN (\partial_reg[7][6] ), .A1 (n_4_0_39), .A2 (n_4_0_7));
NOR2_X1 i_4_0_269 (.ZN (\partial_reg[7][5] ), .A1 (n_4_0_39), .A2 (n_4_0_6));
NOR2_X1 i_4_0_268 (.ZN (\partial_reg[7][4] ), .A1 (n_4_0_39), .A2 (n_4_0_5));
NOR2_X1 i_4_0_267 (.ZN (\partial_reg[7][3] ), .A1 (n_4_0_39), .A2 (n_4_0_4));
NOR2_X1 i_4_0_266 (.ZN (\partial_reg[7][2] ), .A1 (n_4_0_39), .A2 (n_4_0_3));
NOR2_X1 i_4_0_265 (.ZN (\partial_reg[7][1] ), .A1 (n_4_0_39), .A2 (n_4_0_2));
NOR2_X1 i_4_0_264 (.ZN (\partial_reg[7][0] ), .A1 (n_4_0_39), .A2 (n_4_0_1));
INV_X2 i_4_0_263 (.ZN (n_4_0_39), .A (\op2[7] ));
NOR2_X1 i_4_0_262 (.ZN (\partial_reg[6][31] ), .A1 (n_4_0_38), .A2 (n_4_0_32));
NOR2_X1 i_4_0_261 (.ZN (\partial_reg[6][30] ), .A1 (n_4_0_38), .A2 (n_4_0_31));
NOR2_X1 i_4_0_260 (.ZN (\partial_reg[6][29] ), .A1 (n_4_0_38), .A2 (n_4_0_30));
NOR2_X1 i_4_0_259 (.ZN (\partial_reg[6][28] ), .A1 (n_4_0_38), .A2 (n_4_0_29));
NOR2_X1 i_4_0_258 (.ZN (\partial_reg[6][27] ), .A1 (n_4_0_38), .A2 (n_4_0_28));
NOR2_X1 i_4_0_257 (.ZN (\partial_reg[6][26] ), .A1 (n_4_0_38), .A2 (n_4_0_27));
NOR2_X1 i_4_0_256 (.ZN (\partial_reg[6][25] ), .A1 (n_4_0_38), .A2 (n_4_0_26));
NOR2_X1 i_4_0_255 (.ZN (\partial_reg[6][24] ), .A1 (n_4_0_38), .A2 (n_4_0_25));
NOR2_X1 i_4_0_254 (.ZN (\partial_reg[6][23] ), .A1 (n_4_0_38), .A2 (n_4_0_24));
NOR2_X1 i_4_0_253 (.ZN (\partial_reg[6][22] ), .A1 (n_4_0_38), .A2 (n_4_0_23));
NOR2_X1 i_4_0_252 (.ZN (\partial_reg[6][21] ), .A1 (n_4_0_38), .A2 (n_4_0_22));
NOR2_X1 i_4_0_251 (.ZN (\partial_reg[6][20] ), .A1 (n_4_0_38), .A2 (n_4_0_21));
NOR2_X1 i_4_0_250 (.ZN (\partial_reg[6][19] ), .A1 (n_4_0_38), .A2 (n_4_0_20));
NOR2_X1 i_4_0_249 (.ZN (\partial_reg[6][18] ), .A1 (n_4_0_38), .A2 (n_4_0_19));
NOR2_X1 i_4_0_248 (.ZN (\partial_reg[6][17] ), .A1 (n_4_0_38), .A2 (n_4_0_18));
NOR2_X1 i_4_0_247 (.ZN (\partial_reg[6][16] ), .A1 (n_4_0_38), .A2 (n_4_0_17));
NOR2_X1 i_4_0_246 (.ZN (\partial_reg[6][15] ), .A1 (n_4_0_38), .A2 (n_4_0_16));
NOR2_X1 i_4_0_245 (.ZN (\partial_reg[6][14] ), .A1 (n_4_0_38), .A2 (n_4_0_15));
NOR2_X1 i_4_0_244 (.ZN (\partial_reg[6][13] ), .A1 (n_4_0_38), .A2 (n_4_0_14));
NOR2_X1 i_4_0_243 (.ZN (\partial_reg[6][12] ), .A1 (n_4_0_38), .A2 (n_4_0_13));
NOR2_X1 i_4_0_242 (.ZN (\partial_reg[6][11] ), .A1 (n_4_0_38), .A2 (n_4_0_12));
NOR2_X1 i_4_0_241 (.ZN (\partial_reg[6][10] ), .A1 (n_4_0_38), .A2 (n_4_0_11));
NOR2_X1 i_4_0_240 (.ZN (\partial_reg[6][9] ), .A1 (n_4_0_38), .A2 (n_4_0_10));
NOR2_X1 i_4_0_239 (.ZN (\partial_reg[6][8] ), .A1 (n_4_0_38), .A2 (n_4_0_9));
NOR2_X1 i_4_0_238 (.ZN (\partial_reg[6][7] ), .A1 (n_4_0_38), .A2 (n_4_0_8));
NOR2_X1 i_4_0_237 (.ZN (\partial_reg[6][6] ), .A1 (n_4_0_38), .A2 (n_4_0_7));
NOR2_X1 i_4_0_236 (.ZN (\partial_reg[6][5] ), .A1 (n_4_0_38), .A2 (n_4_0_6));
NOR2_X1 i_4_0_235 (.ZN (\partial_reg[6][4] ), .A1 (n_4_0_38), .A2 (n_4_0_5));
NOR2_X1 i_4_0_234 (.ZN (\partial_reg[6][3] ), .A1 (n_4_0_38), .A2 (n_4_0_4));
NOR2_X1 i_4_0_233 (.ZN (\partial_reg[6][2] ), .A1 (n_4_0_38), .A2 (n_4_0_3));
NOR2_X1 i_4_0_232 (.ZN (\partial_reg[6][1] ), .A1 (n_4_0_38), .A2 (n_4_0_2));
NOR2_X1 i_4_0_231 (.ZN (\partial_reg[6][0] ), .A1 (n_4_0_38), .A2 (n_4_0_1));
INV_X2 i_4_0_230 (.ZN (n_4_0_38), .A (\op2[6] ));
NOR2_X1 i_4_0_229 (.ZN (\partial_reg[5][31] ), .A1 (n_4_0_37), .A2 (n_4_0_32));
NOR2_X1 i_4_0_228 (.ZN (\partial_reg[5][30] ), .A1 (n_4_0_37), .A2 (n_4_0_31));
NOR2_X1 i_4_0_227 (.ZN (\partial_reg[5][29] ), .A1 (n_4_0_37), .A2 (n_4_0_30));
NOR2_X1 i_4_0_226 (.ZN (\partial_reg[5][28] ), .A1 (n_4_0_37), .A2 (n_4_0_29));
NOR2_X1 i_4_0_225 (.ZN (\partial_reg[5][27] ), .A1 (n_4_0_37), .A2 (n_4_0_28));
NOR2_X1 i_4_0_224 (.ZN (\partial_reg[5][26] ), .A1 (n_4_0_37), .A2 (n_4_0_27));
NOR2_X1 i_4_0_223 (.ZN (\partial_reg[5][25] ), .A1 (n_4_0_37), .A2 (n_4_0_26));
NOR2_X1 i_4_0_222 (.ZN (\partial_reg[5][24] ), .A1 (n_4_0_37), .A2 (n_4_0_25));
NOR2_X1 i_4_0_221 (.ZN (\partial_reg[5][23] ), .A1 (n_4_0_37), .A2 (n_4_0_24));
NOR2_X1 i_4_0_220 (.ZN (\partial_reg[5][22] ), .A1 (n_4_0_37), .A2 (n_4_0_23));
NOR2_X1 i_4_0_219 (.ZN (\partial_reg[5][21] ), .A1 (n_4_0_37), .A2 (n_4_0_22));
NOR2_X1 i_4_0_218 (.ZN (\partial_reg[5][20] ), .A1 (n_4_0_37), .A2 (n_4_0_21));
NOR2_X1 i_4_0_217 (.ZN (\partial_reg[5][19] ), .A1 (n_4_0_37), .A2 (n_4_0_20));
NOR2_X1 i_4_0_216 (.ZN (\partial_reg[5][18] ), .A1 (n_4_0_37), .A2 (n_4_0_19));
NOR2_X1 i_4_0_215 (.ZN (\partial_reg[5][17] ), .A1 (n_4_0_37), .A2 (n_4_0_18));
NOR2_X1 i_4_0_214 (.ZN (\partial_reg[5][16] ), .A1 (n_4_0_37), .A2 (n_4_0_17));
NOR2_X1 i_4_0_213 (.ZN (\partial_reg[5][15] ), .A1 (n_4_0_37), .A2 (n_4_0_16));
NOR2_X1 i_4_0_212 (.ZN (\partial_reg[5][14] ), .A1 (n_4_0_37), .A2 (n_4_0_15));
NOR2_X1 i_4_0_211 (.ZN (\partial_reg[5][13] ), .A1 (n_4_0_37), .A2 (n_4_0_14));
NOR2_X1 i_4_0_210 (.ZN (\partial_reg[5][12] ), .A1 (n_4_0_37), .A2 (n_4_0_13));
NOR2_X1 i_4_0_209 (.ZN (\partial_reg[5][11] ), .A1 (n_4_0_37), .A2 (n_4_0_12));
NOR2_X1 i_4_0_208 (.ZN (\partial_reg[5][10] ), .A1 (n_4_0_37), .A2 (n_4_0_11));
NOR2_X1 i_4_0_207 (.ZN (\partial_reg[5][9] ), .A1 (n_4_0_37), .A2 (n_4_0_10));
NOR2_X1 i_4_0_206 (.ZN (\partial_reg[5][8] ), .A1 (n_4_0_37), .A2 (n_4_0_9));
NOR2_X1 i_4_0_205 (.ZN (\partial_reg[5][7] ), .A1 (n_4_0_37), .A2 (n_4_0_8));
NOR2_X1 i_4_0_204 (.ZN (\partial_reg[5][6] ), .A1 (n_4_0_37), .A2 (n_4_0_7));
NOR2_X1 i_4_0_203 (.ZN (\partial_reg[5][5] ), .A1 (n_4_0_37), .A2 (n_4_0_6));
NOR2_X1 i_4_0_202 (.ZN (\partial_reg[5][4] ), .A1 (n_4_0_37), .A2 (n_4_0_5));
NOR2_X1 i_4_0_201 (.ZN (\partial_reg[5][3] ), .A1 (n_4_0_37), .A2 (n_4_0_4));
NOR2_X1 i_4_0_200 (.ZN (\partial_reg[5][2] ), .A1 (n_4_0_37), .A2 (n_4_0_3));
NOR2_X1 i_4_0_199 (.ZN (\partial_reg[5][1] ), .A1 (n_4_0_37), .A2 (n_4_0_2));
NOR2_X1 i_4_0_198 (.ZN (\partial_reg[5][0] ), .A1 (n_4_0_37), .A2 (n_4_0_1));
INV_X4 i_4_0_197 (.ZN (n_4_0_37), .A (\op2[5] ));
NOR2_X1 i_4_0_196 (.ZN (\partial_reg[4][31] ), .A1 (n_4_0_36), .A2 (n_4_0_32));
NOR2_X1 i_4_0_195 (.ZN (\partial_reg[4][30] ), .A1 (n_4_0_36), .A2 (n_4_0_31));
NOR2_X1 i_4_0_194 (.ZN (\partial_reg[4][29] ), .A1 (n_4_0_36), .A2 (n_4_0_30));
NOR2_X1 i_4_0_193 (.ZN (\partial_reg[4][28] ), .A1 (n_4_0_36), .A2 (n_4_0_29));
NOR2_X1 i_4_0_192 (.ZN (\partial_reg[4][27] ), .A1 (n_4_0_36), .A2 (n_4_0_28));
NOR2_X1 i_4_0_191 (.ZN (\partial_reg[4][26] ), .A1 (n_4_0_36), .A2 (n_4_0_27));
NOR2_X1 i_4_0_190 (.ZN (\partial_reg[4][25] ), .A1 (n_4_0_36), .A2 (n_4_0_26));
NOR2_X1 i_4_0_189 (.ZN (\partial_reg[4][24] ), .A1 (n_4_0_36), .A2 (n_4_0_25));
NOR2_X1 i_4_0_188 (.ZN (\partial_reg[4][23] ), .A1 (n_4_0_36), .A2 (n_4_0_24));
NOR2_X1 i_4_0_187 (.ZN (\partial_reg[4][22] ), .A1 (n_4_0_36), .A2 (n_4_0_23));
NOR2_X1 i_4_0_186 (.ZN (\partial_reg[4][21] ), .A1 (n_4_0_36), .A2 (n_4_0_22));
NOR2_X1 i_4_0_185 (.ZN (\partial_reg[4][20] ), .A1 (n_4_0_36), .A2 (n_4_0_21));
NOR2_X1 i_4_0_184 (.ZN (\partial_reg[4][19] ), .A1 (n_4_0_36), .A2 (n_4_0_20));
NOR2_X1 i_4_0_183 (.ZN (\partial_reg[4][18] ), .A1 (n_4_0_36), .A2 (n_4_0_19));
NOR2_X1 i_4_0_182 (.ZN (\partial_reg[4][17] ), .A1 (n_4_0_36), .A2 (n_4_0_18));
NOR2_X1 i_4_0_181 (.ZN (\partial_reg[4][16] ), .A1 (n_4_0_36), .A2 (n_4_0_17));
NOR2_X1 i_4_0_180 (.ZN (\partial_reg[4][15] ), .A1 (n_4_0_36), .A2 (n_4_0_16));
NOR2_X1 i_4_0_179 (.ZN (\partial_reg[4][14] ), .A1 (n_4_0_36), .A2 (n_4_0_15));
NOR2_X1 i_4_0_178 (.ZN (\partial_reg[4][13] ), .A1 (n_4_0_36), .A2 (n_4_0_14));
NOR2_X1 i_4_0_177 (.ZN (\partial_reg[4][12] ), .A1 (n_4_0_36), .A2 (n_4_0_13));
NOR2_X1 i_4_0_176 (.ZN (\partial_reg[4][11] ), .A1 (n_4_0_36), .A2 (n_4_0_12));
NOR2_X1 i_4_0_175 (.ZN (\partial_reg[4][10] ), .A1 (n_4_0_36), .A2 (n_4_0_11));
NOR2_X1 i_4_0_174 (.ZN (\partial_reg[4][9] ), .A1 (n_4_0_36), .A2 (n_4_0_10));
NOR2_X1 i_4_0_173 (.ZN (\partial_reg[4][8] ), .A1 (n_4_0_36), .A2 (n_4_0_9));
NOR2_X1 i_4_0_172 (.ZN (\partial_reg[4][7] ), .A1 (n_4_0_36), .A2 (n_4_0_8));
NOR2_X1 i_4_0_171 (.ZN (\partial_reg[4][6] ), .A1 (n_4_0_36), .A2 (n_4_0_7));
NOR2_X1 i_4_0_170 (.ZN (\partial_reg[4][5] ), .A1 (n_4_0_36), .A2 (n_4_0_6));
NOR2_X1 i_4_0_169 (.ZN (\partial_reg[4][4] ), .A1 (n_4_0_36), .A2 (n_4_0_5));
NOR2_X1 i_4_0_168 (.ZN (\partial_reg[4][3] ), .A1 (n_4_0_36), .A2 (n_4_0_4));
NOR2_X1 i_4_0_167 (.ZN (\partial_reg[4][2] ), .A1 (n_4_0_36), .A2 (n_4_0_3));
NOR2_X1 i_4_0_166 (.ZN (\partial_reg[4][1] ), .A1 (n_4_0_36), .A2 (n_4_0_2));
NOR2_X1 i_4_0_165 (.ZN (\partial_reg[4][0] ), .A1 (n_4_0_36), .A2 (n_4_0_1));
INV_X4 i_4_0_164 (.ZN (n_4_0_36), .A (\op2[4] ));
NOR2_X1 i_4_0_163 (.ZN (\partial_reg[3][31] ), .A1 (n_4_0_35), .A2 (n_4_0_32));
NOR2_X1 i_4_0_162 (.ZN (\partial_reg[3][30] ), .A1 (n_4_0_35), .A2 (n_4_0_31));
NOR2_X1 i_4_0_161 (.ZN (\partial_reg[3][29] ), .A1 (n_4_0_35), .A2 (n_4_0_30));
NOR2_X1 i_4_0_160 (.ZN (\partial_reg[3][28] ), .A1 (n_4_0_35), .A2 (n_4_0_29));
NOR2_X1 i_4_0_159 (.ZN (\partial_reg[3][27] ), .A1 (n_4_0_35), .A2 (n_4_0_28));
NOR2_X1 i_4_0_158 (.ZN (\partial_reg[3][26] ), .A1 (n_4_0_35), .A2 (n_4_0_27));
NOR2_X1 i_4_0_157 (.ZN (\partial_reg[3][25] ), .A1 (n_4_0_35), .A2 (n_4_0_26));
NOR2_X1 i_4_0_156 (.ZN (\partial_reg[3][24] ), .A1 (n_4_0_35), .A2 (n_4_0_25));
NOR2_X1 i_4_0_155 (.ZN (\partial_reg[3][23] ), .A1 (n_4_0_35), .A2 (n_4_0_24));
NOR2_X1 i_4_0_154 (.ZN (\partial_reg[3][22] ), .A1 (n_4_0_35), .A2 (n_4_0_23));
NOR2_X1 i_4_0_153 (.ZN (\partial_reg[3][21] ), .A1 (n_4_0_35), .A2 (n_4_0_22));
NOR2_X1 i_4_0_152 (.ZN (\partial_reg[3][20] ), .A1 (n_4_0_35), .A2 (n_4_0_21));
NOR2_X1 i_4_0_151 (.ZN (\partial_reg[3][19] ), .A1 (n_4_0_35), .A2 (n_4_0_20));
NOR2_X1 i_4_0_150 (.ZN (\partial_reg[3][18] ), .A1 (n_4_0_35), .A2 (n_4_0_19));
NOR2_X1 i_4_0_149 (.ZN (\partial_reg[3][17] ), .A1 (n_4_0_35), .A2 (n_4_0_18));
NOR2_X1 i_4_0_148 (.ZN (\partial_reg[3][16] ), .A1 (n_4_0_35), .A2 (n_4_0_17));
NOR2_X1 i_4_0_147 (.ZN (\partial_reg[3][15] ), .A1 (n_4_0_35), .A2 (n_4_0_16));
NOR2_X1 i_4_0_146 (.ZN (\partial_reg[3][14] ), .A1 (n_4_0_35), .A2 (n_4_0_15));
NOR2_X1 i_4_0_145 (.ZN (\partial_reg[3][13] ), .A1 (n_4_0_35), .A2 (n_4_0_14));
NOR2_X1 i_4_0_144 (.ZN (\partial_reg[3][12] ), .A1 (n_4_0_35), .A2 (n_4_0_13));
NOR2_X1 i_4_0_143 (.ZN (\partial_reg[3][11] ), .A1 (n_4_0_35), .A2 (n_4_0_12));
NOR2_X1 i_4_0_142 (.ZN (\partial_reg[3][10] ), .A1 (n_4_0_35), .A2 (n_4_0_11));
NOR2_X1 i_4_0_141 (.ZN (\partial_reg[3][9] ), .A1 (n_4_0_35), .A2 (n_4_0_10));
NOR2_X1 i_4_0_140 (.ZN (\partial_reg[3][8] ), .A1 (n_4_0_35), .A2 (n_4_0_9));
NOR2_X1 i_4_0_139 (.ZN (\partial_reg[3][7] ), .A1 (n_4_0_35), .A2 (n_4_0_8));
NOR2_X1 i_4_0_138 (.ZN (\partial_reg[3][6] ), .A1 (n_4_0_35), .A2 (n_4_0_7));
NOR2_X1 i_4_0_137 (.ZN (\partial_reg[3][5] ), .A1 (n_4_0_35), .A2 (n_4_0_6));
NOR2_X1 i_4_0_136 (.ZN (\partial_reg[3][4] ), .A1 (n_4_0_35), .A2 (n_4_0_5));
NOR2_X1 i_4_0_135 (.ZN (\partial_reg[3][3] ), .A1 (n_4_0_35), .A2 (n_4_0_4));
NOR2_X1 i_4_0_134 (.ZN (\partial_reg[3][2] ), .A1 (n_4_0_35), .A2 (n_4_0_3));
NOR2_X1 i_4_0_133 (.ZN (\partial_reg[3][1] ), .A1 (n_4_0_35), .A2 (n_4_0_2));
NOR2_X1 i_4_0_132 (.ZN (\partial_reg[3][0] ), .A1 (n_4_0_35), .A2 (n_4_0_1));
INV_X2 i_4_0_131 (.ZN (n_4_0_35), .A (\op2[3] ));
NOR2_X1 i_4_0_130 (.ZN (\partial_reg[2][31] ), .A1 (n_4_0_34), .A2 (n_4_0_32));
NOR2_X1 i_4_0_127 (.ZN (\partial_reg[2][28] ), .A1 (n_4_0_34), .A2 (n_4_0_29));
NOR2_X1 i_4_0_126 (.ZN (\partial_reg[2][27] ), .A1 (n_4_0_34), .A2 (n_4_0_28));
NOR2_X1 i_4_0_125 (.ZN (\partial_reg[2][26] ), .A1 (n_4_0_34), .A2 (n_4_0_27));
NOR2_X1 i_4_0_124 (.ZN (\partial_reg[2][25] ), .A1 (n_4_0_34), .A2 (n_4_0_26));
NOR2_X1 i_4_0_123 (.ZN (\partial_reg[2][24] ), .A1 (n_4_0_34), .A2 (n_4_0_25));
NOR2_X1 i_4_0_122 (.ZN (\partial_reg[2][23] ), .A1 (n_4_0_34), .A2 (n_4_0_24));
NOR2_X1 i_4_0_121 (.ZN (\partial_reg[2][22] ), .A1 (n_4_0_34), .A2 (n_4_0_23));
NOR2_X1 i_4_0_120 (.ZN (\partial_reg[2][21] ), .A1 (n_4_0_34), .A2 (n_4_0_22));
NOR2_X2 i_4_0_119 (.ZN (\partial_reg[2][20] ), .A1 (n_4_0_34), .A2 (n_4_0_21));
NOR2_X2 i_4_0_118 (.ZN (\partial_reg[2][19] ), .A1 (n_4_0_34), .A2 (n_4_0_20));
NOR2_X1 i_4_0_117 (.ZN (\partial_reg[2][18] ), .A1 (n_4_0_34), .A2 (n_4_0_19));
NOR2_X1 i_4_0_116 (.ZN (\partial_reg[2][17] ), .A1 (n_4_0_34), .A2 (n_4_0_18));
NOR2_X1 i_4_0_115 (.ZN (\partial_reg[2][16] ), .A1 (n_4_0_34), .A2 (n_4_0_17));
NOR2_X1 i_4_0_114 (.ZN (\partial_reg[2][15] ), .A1 (n_4_0_34), .A2 (n_4_0_16));
NOR2_X1 i_4_0_113 (.ZN (\partial_reg[2][14] ), .A1 (n_4_0_34), .A2 (n_4_0_15));
NOR2_X1 i_4_0_112 (.ZN (\partial_reg[2][13] ), .A1 (n_4_0_34), .A2 (n_4_0_14));
NOR2_X1 i_4_0_111 (.ZN (\partial_reg[2][12] ), .A1 (n_4_0_34), .A2 (n_4_0_13));
NOR2_X1 i_4_0_110 (.ZN (\partial_reg[2][11] ), .A1 (n_4_0_34), .A2 (n_4_0_12));
NOR2_X1 i_4_0_109 (.ZN (\partial_reg[2][10] ), .A1 (n_4_0_34), .A2 (n_4_0_11));
NOR2_X1 i_4_0_108 (.ZN (\partial_reg[2][9] ), .A1 (n_4_0_34), .A2 (n_4_0_10));
NOR2_X1 i_4_0_107 (.ZN (\partial_reg[2][8] ), .A1 (n_4_0_34), .A2 (n_4_0_9));
NOR2_X1 i_4_0_106 (.ZN (\partial_reg[2][7] ), .A1 (n_4_0_34), .A2 (n_4_0_8));
NOR2_X1 i_4_0_105 (.ZN (\partial_reg[2][6] ), .A1 (n_4_0_34), .A2 (n_4_0_7));
NOR2_X1 i_4_0_104 (.ZN (\partial_reg[2][5] ), .A1 (n_4_0_34), .A2 (n_4_0_6));
NOR2_X1 i_4_0_103 (.ZN (\partial_reg[2][4] ), .A1 (n_4_0_34), .A2 (n_4_0_5));
NOR2_X1 i_4_0_102 (.ZN (\partial_reg[2][3] ), .A1 (n_4_0_34), .A2 (n_4_0_4));
NOR2_X1 i_4_0_101 (.ZN (\partial_reg[2][2] ), .A1 (n_4_0_34), .A2 (n_4_0_3));
NOR2_X1 i_4_0_100 (.ZN (\partial_reg[2][1] ), .A1 (n_4_0_34), .A2 (n_4_0_2));
NOR2_X1 i_4_0_99 (.ZN (\partial_reg[2][0] ), .A1 (n_4_0_34), .A2 (n_4_0_1));
NOR2_X1 i_4_0_95 (.ZN (\partial_reg[1][29] ), .A1 (n_4_0_33), .A2 (n_4_0_30));
NOR2_X1 i_4_0_94 (.ZN (\partial_reg[1][28] ), .A1 (n_4_0_33), .A2 (n_4_0_29));
NOR2_X1 i_4_0_93 (.ZN (\partial_reg[1][27] ), .A1 (n_4_0_33), .A2 (n_4_0_28));
NOR2_X1 i_4_0_92 (.ZN (\partial_reg[1][26] ), .A1 (n_4_0_33), .A2 (n_4_0_27));
NOR2_X1 i_4_0_91 (.ZN (\partial_reg[1][25] ), .A1 (n_4_0_33), .A2 (n_4_0_26));
NOR2_X1 i_4_0_90 (.ZN (\partial_reg[1][24] ), .A1 (n_4_0_33), .A2 (n_4_0_25));
NOR2_X1 i_4_0_89 (.ZN (\partial_reg[1][23] ), .A1 (n_4_0_33), .A2 (n_4_0_24));
NOR2_X1 i_4_0_88 (.ZN (\partial_reg[1][22] ), .A1 (n_4_0_33), .A2 (n_4_0_23));
NOR2_X1 i_4_0_87 (.ZN (\partial_reg[1][21] ), .A1 (n_4_0_33), .A2 (n_4_0_22));
NOR2_X1 i_4_0_86 (.ZN (\partial_reg[1][20] ), .A1 (n_4_0_33), .A2 (n_4_0_21));
NOR2_X1 i_4_0_85 (.ZN (\partial_reg[1][19] ), .A1 (n_4_0_33), .A2 (n_4_0_20));
NOR2_X1 i_4_0_84 (.ZN (\partial_reg[1][18] ), .A1 (n_4_0_33), .A2 (n_4_0_19));
NOR2_X1 i_4_0_83 (.ZN (\partial_reg[1][17] ), .A1 (n_4_0_33), .A2 (n_4_0_18));
NOR2_X1 i_4_0_82 (.ZN (\partial_reg[1][16] ), .A1 (n_4_0_33), .A2 (n_4_0_17));
NOR2_X1 i_4_0_81 (.ZN (\partial_reg[1][15] ), .A1 (n_4_0_33), .A2 (n_4_0_16));
NOR2_X1 i_4_0_80 (.ZN (\partial_reg[1][14] ), .A1 (n_4_0_33), .A2 (n_4_0_15));
NOR2_X1 i_4_0_79 (.ZN (\partial_reg[1][13] ), .A1 (n_4_0_33), .A2 (n_4_0_14));
NOR2_X1 i_4_0_78 (.ZN (\partial_reg[1][12] ), .A1 (n_4_0_33), .A2 (n_4_0_13));
NOR2_X1 i_4_0_77 (.ZN (\partial_reg[1][11] ), .A1 (n_4_0_33), .A2 (n_4_0_12));
NOR2_X1 i_4_0_76 (.ZN (\partial_reg[1][10] ), .A1 (n_4_0_33), .A2 (n_4_0_11));
NOR2_X1 i_4_0_75 (.ZN (\partial_reg[1][9] ), .A1 (n_4_0_33), .A2 (n_4_0_10));
NOR2_X1 i_4_0_74 (.ZN (\partial_reg[1][8] ), .A1 (n_4_0_33), .A2 (n_4_0_9));
NOR2_X1 i_4_0_73 (.ZN (\partial_reg[1][7] ), .A1 (n_4_0_33), .A2 (n_4_0_8));
NOR2_X1 i_4_0_72 (.ZN (\partial_reg[1][6] ), .A1 (n_4_0_33), .A2 (n_4_0_7));
NOR2_X1 i_4_0_71 (.ZN (\partial_reg[1][5] ), .A1 (n_4_0_33), .A2 (n_4_0_6));
NOR2_X1 i_4_0_70 (.ZN (\partial_reg[1][4] ), .A1 (n_4_0_33), .A2 (n_4_0_5));
NOR2_X1 i_4_0_69 (.ZN (\partial_reg[1][3] ), .A1 (n_4_0_33), .A2 (n_4_0_4));
NOR2_X1 i_4_0_68 (.ZN (\partial_reg[1][2] ), .A1 (n_4_0_33), .A2 (n_4_0_3));
NOR2_X1 i_4_0_67 (.ZN (\partial_reg[1][1] ), .A1 (n_4_0_33), .A2 (n_4_0_2));
NOR2_X1 i_4_0_66 (.ZN (\partial_reg[1][0] ), .A1 (n_4_0_33), .A2 (n_4_0_1));
NOR2_X1 i_4_0_62 (.ZN (\partial_reg[0][30] ), .A1 (n_4_0_0), .A2 (n_4_0_31));
NOR2_X1 i_4_0_60 (.ZN (\partial_reg[0][29] ), .A1 (n_4_0_0), .A2 (n_4_0_30));
NOR2_X2 i_4_0_58 (.ZN (\partial_reg[0][28] ), .A1 (n_4_0_0), .A2 (n_4_0_29));
INV_X2 i_4_0_57 (.ZN (n_4_0_29), .A (\op1[28] ));
NOR2_X1 i_4_0_56 (.ZN (\partial_reg[0][27] ), .A1 (n_4_0_0), .A2 (n_4_0_28));
INV_X2 i_4_0_55 (.ZN (n_4_0_28), .A (\op1[27] ));
NOR2_X2 i_4_0_54 (.ZN (\partial_reg[0][26] ), .A1 (n_4_0_0), .A2 (n_4_0_27));
INV_X8 i_4_0_53 (.ZN (n_4_0_27), .A (\op1[26] ));
NOR2_X2 i_4_0_52 (.ZN (\partial_reg[0][25] ), .A1 (n_4_0_0), .A2 (n_4_0_26));
INV_X4 i_4_0_51 (.ZN (n_4_0_26), .A (\op1[25] ));
NOR2_X2 i_4_0_50 (.ZN (\partial_reg[0][24] ), .A1 (n_4_0_0), .A2 (n_4_0_25));
INV_X8 i_4_0_49 (.ZN (n_4_0_25), .A (\op1[24] ));
NOR2_X1 i_4_0_48 (.ZN (\partial_reg[0][23] ), .A1 (n_4_0_0), .A2 (n_4_0_24));
INV_X4 i_4_0_47 (.ZN (n_4_0_24), .A (\op1[23] ));
NOR2_X2 i_4_0_46 (.ZN (\partial_reg[0][22] ), .A1 (n_4_0_0), .A2 (n_4_0_23));
INV_X4 i_4_0_45 (.ZN (n_4_0_23), .A (\op1[22] ));
NOR2_X1 i_4_0_44 (.ZN (\partial_reg[0][21] ), .A1 (n_4_0_0), .A2 (n_4_0_22));
INV_X4 i_4_0_43 (.ZN (n_4_0_22), .A (\op1[21] ));
NOR2_X1 i_4_0_42 (.ZN (\partial_reg[0][20] ), .A1 (n_4_0_0), .A2 (n_4_0_21));
INV_X4 i_4_0_41 (.ZN (n_4_0_21), .A (\op1[20] ));
NOR2_X1 i_4_0_40 (.ZN (\partial_reg[0][19] ), .A1 (n_4_0_0), .A2 (n_4_0_20));
INV_X4 i_4_0_39 (.ZN (n_4_0_20), .A (\op1[19] ));
NOR2_X1 i_4_0_38 (.ZN (\partial_reg[0][18] ), .A1 (n_4_0_0), .A2 (n_4_0_19));
INV_X2 i_4_0_37 (.ZN (n_4_0_19), .A (\op1[18] ));
NOR2_X1 i_4_0_36 (.ZN (\partial_reg[0][17] ), .A1 (n_4_0_0), .A2 (n_4_0_18));
INV_X2 i_4_0_35 (.ZN (n_4_0_18), .A (\op1[17] ));
NOR2_X1 i_4_0_34 (.ZN (\partial_reg[0][16] ), .A1 (n_4_0_0), .A2 (n_4_0_17));
INV_X2 i_4_0_33 (.ZN (n_4_0_17), .A (\op1[16] ));
NOR2_X1 i_4_0_32 (.ZN (\partial_reg[0][15] ), .A1 (n_4_0_0), .A2 (n_4_0_16));
INV_X2 i_4_0_31 (.ZN (n_4_0_16), .A (\op1[15] ));
NOR2_X1 i_4_0_30 (.ZN (\partial_reg[0][14] ), .A1 (n_4_0_0), .A2 (n_4_0_15));
INV_X2 i_4_0_29 (.ZN (n_4_0_15), .A (\op1[14] ));
NOR2_X1 i_4_0_28 (.ZN (\partial_reg[0][13] ), .A1 (n_4_0_0), .A2 (n_4_0_14));
INV_X2 i_4_0_27 (.ZN (n_4_0_14), .A (\op1[13] ));
NOR2_X1 i_4_0_26 (.ZN (\partial_reg[0][12] ), .A1 (n_4_0_0), .A2 (n_4_0_13));
INV_X2 i_4_0_25 (.ZN (n_4_0_13), .A (\op1[12] ));
NOR2_X1 i_4_0_24 (.ZN (\partial_reg[0][11] ), .A1 (n_4_0_0), .A2 (n_4_0_12));
INV_X2 i_4_0_23 (.ZN (n_4_0_12), .A (\op1[11] ));
NOR2_X1 i_4_0_22 (.ZN (\partial_reg[0][10] ), .A1 (n_4_0_0), .A2 (n_4_0_11));
INV_X2 i_4_0_21 (.ZN (n_4_0_11), .A (\op1[10] ));
NOR2_X1 i_4_0_20 (.ZN (\partial_reg[0][9] ), .A1 (n_4_0_0), .A2 (n_4_0_10));
INV_X2 i_4_0_19 (.ZN (n_4_0_10), .A (\op1[9] ));
NOR2_X1 i_4_0_18 (.ZN (\partial_reg[0][8] ), .A1 (n_4_0_0), .A2 (n_4_0_9));
INV_X2 i_4_0_17 (.ZN (n_4_0_9), .A (\op1[8] ));
NOR2_X1 i_4_0_16 (.ZN (\partial_reg[0][7] ), .A1 (n_4_0_0), .A2 (n_4_0_8));
INV_X2 i_4_0_15 (.ZN (n_4_0_8), .A (\op1[7] ));
NOR2_X1 i_4_0_14 (.ZN (\partial_reg[0][6] ), .A1 (n_4_0_0), .A2 (n_4_0_7));
INV_X2 i_4_0_13 (.ZN (n_4_0_7), .A (\op1[6] ));
NOR2_X1 i_4_0_12 (.ZN (\partial_reg[0][5] ), .A1 (n_4_0_0), .A2 (n_4_0_6));
INV_X2 i_4_0_11 (.ZN (n_4_0_6), .A (\op1[5] ));
NOR2_X1 i_4_0_10 (.ZN (\partial_reg[0][4] ), .A1 (n_4_0_0), .A2 (n_4_0_5));
INV_X2 i_4_0_9 (.ZN (n_4_0_5), .A (\op1[4] ));
NOR2_X1 i_4_0_8 (.ZN (\partial_reg[0][3] ), .A1 (n_4_0_0), .A2 (n_4_0_4));
INV_X2 i_4_0_7 (.ZN (n_4_0_4), .A (\op1[3] ));
NOR2_X1 i_4_0_6 (.ZN (\partial_reg[0][2] ), .A1 (n_4_0_0), .A2 (n_4_0_3));
INV_X2 i_4_0_5 (.ZN (n_4_0_3), .A (\op1[2] ));
NOR2_X1 i_4_0_4 (.ZN (\partial_reg[0][1] ), .A1 (n_4_0_0), .A2 (n_4_0_2));
INV_X2 i_4_0_3 (.ZN (n_4_0_2), .A (\op1[1] ));
NOR2_X1 i_4_0_2 (.ZN (out[0]), .A1 (n_4_0_0), .A2 (n_4_0_1));
INV_X2 i_4_0_1 (.ZN (n_4_0_1), .A (a[0]));
adderPlus final (.cout (n_28), .sum ({n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
    n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, 
    n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29}), .a ({\partial_reg[31][31] , 
    \s1[29][31] , \s1[29][30] , \s1[29][29] , \s1[29][28] , \s1[29][27] , \s1[29][26] , 
    \s1[29][25] , \s1[29][24] , \s1[29][23] , \s1[29][22] , \s1[29][21] , \s1[29][20] , 
    \s1[29][19] , \s1[29][18] , \s1[29][17] , \s1[29][16] , \s1[29][15] , \s1[29][14] , 
    \s1[29][13] , \s1[29][12] , \s1[29][11] , \s1[29][10] , \s1[29][9] , \s1[29][8] , 
    \s1[29][7] , \s1[29][6] , \s1[29][5] , \s1[29][4] , \s1[29][3] , \s1[29][2] , 
    \s1[29][1] }), .b ({\c1[29][31] , \c1[29][30] , \c1[29][29] , \c1[29][28] , \c1[29][27] , 
    \c1[29][26] , \c1[29][25] , \c1[29][24] , \c1[29][23] , \c1[29][22] , \c1[29][21] , 
    \c1[29][20] , \c1[29][19] , \c1[29][18] , \c1[29][17] , \c1[29][16] , \c1[29][15] , 
    \c1[29][14] , \c1[29][13] , \c1[29][12] , \c1[29][11] , \c1[29][10] , \c1[29][9] , 
    \c1[29][8] , \c1[29][7] , \c1[29][6] , \c1[29][5] , \c1[29][4] , \c1[29][3] , 
    \c1[29][2] , \c1[29][1] , \c1[29][0] }));
PartialAdder__0_47 genblk1_29_p2 (.c1 ({\c1[29][31] , \c1[29][30] , \c1[29][29] , 
    \c1[29][28] , \c1[29][27] , \c1[29][26] , \c1[29][25] , \c1[29][24] , \c1[29][23] , 
    \c1[29][22] , \c1[29][21] , \c1[29][20] , \c1[29][19] , \c1[29][18] , \c1[29][17] , 
    \c1[29][16] , \c1[29][15] , \c1[29][14] , \c1[29][13] , \c1[29][12] , \c1[29][11] , 
    \c1[29][10] , \c1[29][9] , \c1[29][8] , \c1[29][7] , \c1[29][6] , \c1[29][5] , 
    \c1[29][4] , \c1[29][3] , \c1[29][2] , \c1[29][1] , \c1[29][0] }), .s1 ({uc_86, 
    \s1[29][31] , \s1[29][30] , \s1[29][29] , \s1[29][28] , \s1[29][27] , \s1[29][26] , 
    \s1[29][25] , \s1[29][24] , \s1[29][23] , \s1[29][22] , \s1[29][21] , \s1[29][20] , 
    \s1[29][19] , \s1[29][18] , \s1[29][17] , \s1[29][16] , \s1[29][15] , \s1[29][14] , 
    \s1[29][13] , \s1[29][12] , \s1[29][11] , \s1[29][10] , \s1[29][9] , \s1[29][8] , 
    \s1[29][7] , \s1[29][6] , \s1[29][5] , \s1[29][4] , \s1[29][3] , \s1[29][2] , 
    \s1[29][1] , \s1[29][0] }), .a ({\partial_reg[30][31] , n_39_863, n_39_831, n_39_799, 
    n_39_767, n_39_735, n_39_703, n_39_671, n_39_639, n_39_607, n_39_575, n_39_543, 
    n_39_511, n_39_479, n_39_447, n_39_415, n_39_383, n_39_351, n_39_319, n_39_287, 
    n_39_255, n_39_223, n_39_191, n_39_159, n_39_127, n_39_95, n_39_63, n_39_31, 
    n_39_867, n_39_866, n_39_865, n_39_864, uc_84}), .b ({\c1[28][31] , \c1[28][30] , 
    \c1[28][29] , \c1[28][28] , \c1[28][27] , \c1[28][26] , \c1[28][25] , \c1[28][24] , 
    \c1[28][23] , \c1[28][22] , \c1[28][21] , \c1[28][20] , \c1[28][19] , \c1[28][18] , 
    \c1[28][17] , \c1[28][16] , \c1[28][15] , \c1[28][14] , \c1[28][13] , \c1[28][12] , 
    \c1[28][11] , \c1[28][10] , \c1[28][9] , \c1[28][8] , \c1[28][7] , \c1[28][6] , 
    \c1[28][5] , \c1[28][4] , \c1[28][3] , \c1[28][2] , \c1[28][1] , \c1[28][0] })
    , .c ({uc_85, \partial_reg[31][30] , \partial_reg[31][29] , \partial_reg[31][28] , 
    \partial_reg[31][27] , \partial_reg[31][26] , \partial_reg[31][25] , \partial_reg[31][24] , 
    \partial_reg[31][23] , \partial_reg[31][22] , \partial_reg[31][21] , \partial_reg[31][20] , 
    \partial_reg[31][19] , \partial_reg[31][18] , \partial_reg[31][17] , \partial_reg[31][16] , 
    \partial_reg[31][15] , \partial_reg[31][14] , \partial_reg[31][13] , \partial_reg[31][12] , 
    \partial_reg[31][11] , \partial_reg[31][10] , \partial_reg[31][9] , \partial_reg[31][8] , 
    \partial_reg[31][7] , \partial_reg[31][6] , \partial_reg[31][5] , \partial_reg[31][4] , 
    \partial_reg[31][3] , \partial_reg[31][2] , \partial_reg[31][1] , \partial_reg[31][0] }));
PartialAdder__1_2805 genblk1_28_p2 (.c1 ({\c1[28][31] , \c1[28][30] , \c1[28][29] , 
    \c1[28][28] , \c1[28][27] , \c1[28][26] , \c1[28][25] , \c1[28][24] , \c1[28][23] , 
    \c1[28][22] , \c1[28][21] , \c1[28][20] , \c1[28][19] , \c1[28][18] , \c1[28][17] , 
    \c1[28][16] , \c1[28][15] , \c1[28][14] , \c1[28][13] , \c1[28][12] , \c1[28][11] , 
    \c1[28][10] , \c1[28][9] , \c1[28][8] , \c1[28][7] , \c1[28][6] , \c1[28][5] , 
    \c1[28][4] , \c1[28][3] , \c1[28][2] , \c1[28][1] , \c1[28][0] }), .s1 ({uc_83, 
    n_39_863, n_39_831, n_39_799, n_39_767, n_39_735, n_39_703, n_39_671, n_39_639, 
    n_39_607, n_39_575, n_39_543, n_39_511, n_39_479, n_39_447, n_39_415, n_39_383, 
    n_39_351, n_39_319, n_39_287, n_39_255, n_39_223, n_39_191, n_39_159, n_39_127, 
    n_39_95, n_39_63, n_39_31, n_39_867, n_39_866, n_39_865, n_39_864, n_27}), .a ({
    \partial_reg[29][31] , n_39_862, n_39_861, n_39_860, n_39_859, n_39_858, n_39_857, 
    n_39_856, n_39_855, n_39_854, n_39_853, n_39_852, n_39_851, n_39_850, n_39_849, 
    n_39_848, n_39_847, n_39_846, n_39_845, n_39_844, n_39_843, n_39_842, n_39_841, 
    n_39_840, n_39_839, n_39_838, n_39_837, n_39_836, n_39_835, n_39_834, n_39_833, 
    n_39_832, uc_81}), .b ({\c1[27][31] , \c1[27][30] , \c1[27][29] , \c1[27][28] , 
    \c1[27][27] , \c1[27][26] , \c1[27][25] , \c1[27][24] , \c1[27][23] , \c1[27][22] , 
    \c1[27][21] , \c1[27][20] , \c1[27][19] , \c1[27][18] , \c1[27][17] , \c1[27][16] , 
    \c1[27][15] , \c1[27][14] , \c1[27][13] , \c1[27][12] , \c1[27][11] , \c1[27][10] , 
    \c1[27][9] , \c1[27][8] , \c1[27][7] , \c1[27][6] , \c1[27][5] , \c1[27][4] , 
    \c1[27][3] , \c1[27][2] , \c1[27][1] , \c1[27][0] }), .c ({uc_82, \partial_reg[30][30] , 
    \partial_reg[30][29] , \partial_reg[30][28] , \partial_reg[30][27] , \partial_reg[30][26] , 
    \partial_reg[30][25] , \partial_reg[30][24] , \partial_reg[30][23] , \partial_reg[30][22] , 
    \partial_reg[30][21] , \partial_reg[30][20] , \partial_reg[30][19] , \partial_reg[30][18] , 
    \partial_reg[30][17] , \partial_reg[30][16] , \partial_reg[30][15] , \partial_reg[30][14] , 
    \partial_reg[30][13] , \partial_reg[30][12] , \partial_reg[30][11] , \partial_reg[30][10] , 
    \partial_reg[30][9] , \partial_reg[30][8] , \partial_reg[30][7] , \partial_reg[30][6] , 
    \partial_reg[30][5] , \partial_reg[30][4] , \partial_reg[30][3] , \partial_reg[30][2] , 
    \partial_reg[30][1] , \partial_reg[30][0] }));
PartialAdder__1_2708 genblk1_27_p2 (.c1 ({\c1[27][31] , \c1[27][30] , \c1[27][29] , 
    \c1[27][28] , \c1[27][27] , \c1[27][26] , \c1[27][25] , \c1[27][24] , \c1[27][23] , 
    \c1[27][22] , \c1[27][21] , \c1[27][20] , \c1[27][19] , \c1[27][18] , \c1[27][17] , 
    \c1[27][16] , \c1[27][15] , \c1[27][14] , \c1[27][13] , \c1[27][12] , \c1[27][11] , 
    \c1[27][10] , \c1[27][9] , \c1[27][8] , \c1[27][7] , \c1[27][6] , \c1[27][5] , 
    \c1[27][4] , \c1[27][3] , \c1[27][2] , \c1[27][1] , \c1[27][0] }), .s1 ({uc_80, 
    n_39_862, n_39_861, n_39_860, n_39_859, n_39_858, n_39_857, n_39_856, n_39_855, 
    n_39_854, n_39_853, n_39_852, n_39_851, n_39_850, n_39_849, n_39_848, n_39_847, 
    n_39_846, n_39_845, n_39_844, n_39_843, n_39_842, n_39_841, n_39_840, n_39_839, 
    n_39_838, n_39_837, n_39_836, n_39_835, n_39_834, n_39_833, n_39_832, n_26}), .a ({
    \partial_reg[28][31] , n_39_830, n_39_829, n_39_828, n_39_827, n_39_826, n_39_825, 
    n_39_824, n_39_823, n_39_822, n_39_821, n_39_820, n_39_819, n_39_818, n_39_817, 
    n_39_816, n_39_815, n_39_814, n_39_813, n_39_812, n_39_811, n_39_810, n_39_809, 
    n_39_808, n_39_807, n_39_806, n_39_805, n_39_804, n_39_803, n_39_802, n_39_801, 
    n_39_800, uc_78}), .b ({\c1[26][31] , \c1[26][30] , \c1[26][29] , \c1[26][28] , 
    \c1[26][27] , \c1[26][26] , \c1[26][25] , \c1[26][24] , \c1[26][23] , \c1[26][22] , 
    \c1[26][21] , \c1[26][20] , \c1[26][19] , \c1[26][18] , \c1[26][17] , \c1[26][16] , 
    \c1[26][15] , \c1[26][14] , \c1[26][13] , \c1[26][12] , \c1[26][11] , \c1[26][10] , 
    \c1[26][9] , \c1[26][8] , \c1[26][7] , \c1[26][6] , \c1[26][5] , \c1[26][4] , 
    \c1[26][3] , \c1[26][2] , \c1[26][1] , \c1[26][0] }), .c ({uc_79, \partial_reg[29][30] , 
    \partial_reg[29][29] , \partial_reg[29][28] , \partial_reg[29][27] , \partial_reg[29][26] , 
    \partial_reg[29][25] , \partial_reg[29][24] , \partial_reg[29][23] , \partial_reg[29][22] , 
    \partial_reg[29][21] , \partial_reg[29][20] , \partial_reg[29][19] , \partial_reg[29][18] , 
    \partial_reg[29][17] , \partial_reg[29][16] , \partial_reg[29][15] , \partial_reg[29][14] , 
    \partial_reg[29][13] , \partial_reg[29][12] , \partial_reg[29][11] , \partial_reg[29][10] , 
    \partial_reg[29][9] , \partial_reg[29][8] , \partial_reg[29][7] , \partial_reg[29][6] , 
    \partial_reg[29][5] , \partial_reg[29][4] , \partial_reg[29][3] , \partial_reg[29][2] , 
    \partial_reg[29][1] , \partial_reg[29][0] }));
PartialAdder__1_2611 genblk1_26_p2 (.c1 ({\c1[26][31] , \c1[26][30] , \c1[26][29] , 
    \c1[26][28] , \c1[26][27] , \c1[26][26] , \c1[26][25] , \c1[26][24] , \c1[26][23] , 
    \c1[26][22] , \c1[26][21] , \c1[26][20] , \c1[26][19] , \c1[26][18] , \c1[26][17] , 
    \c1[26][16] , \c1[26][15] , \c1[26][14] , \c1[26][13] , \c1[26][12] , \c1[26][11] , 
    \c1[26][10] , \c1[26][9] , \c1[26][8] , \c1[26][7] , \c1[26][6] , \c1[26][5] , 
    \c1[26][4] , \c1[26][3] , \c1[26][2] , \c1[26][1] , \c1[26][0] }), .s1 ({uc_77, 
    n_39_830, n_39_829, n_39_828, n_39_827, n_39_826, n_39_825, n_39_824, n_39_823, 
    n_39_822, n_39_821, n_39_820, n_39_819, n_39_818, n_39_817, n_39_816, n_39_815, 
    n_39_814, n_39_813, n_39_812, n_39_811, n_39_810, n_39_809, n_39_808, n_39_807, 
    n_39_806, n_39_805, n_39_804, n_39_803, n_39_802, n_39_801, n_39_800, n_25}), .a ({
    \partial_reg[27][31] , n_39_798, n_39_797, n_39_796, n_39_795, n_39_794, n_39_793, 
    n_39_792, n_39_791, n_39_790, n_39_789, n_39_788, n_39_787, n_39_786, n_39_785, 
    n_39_784, n_39_783, n_39_782, n_39_781, n_39_780, n_39_779, n_39_778, n_39_777, 
    n_39_776, n_39_775, n_39_774, n_39_773, n_39_772, n_39_771, n_39_770, n_39_769, 
    n_39_768, uc_75}), .b ({\c1[25][31] , \c1[25][30] , \c1[25][29] , \c1[25][28] , 
    \c1[25][27] , \c1[25][26] , \c1[25][25] , \c1[25][24] , \c1[25][23] , \c1[25][22] , 
    \c1[25][21] , \c1[25][20] , \c1[25][19] , \c1[25][18] , \c1[25][17] , \c1[25][16] , 
    \c1[25][15] , \c1[25][14] , \c1[25][13] , \c1[25][12] , \c1[25][11] , \c1[25][10] , 
    \c1[25][9] , \c1[25][8] , \c1[25][7] , \c1[25][6] , \c1[25][5] , \c1[25][4] , 
    \c1[25][3] , \c1[25][2] , \c1[25][1] , \c1[25][0] }), .c ({uc_76, \partial_reg[28][30] , 
    \partial_reg[28][29] , \partial_reg[28][28] , \partial_reg[28][27] , \partial_reg[28][26] , 
    \partial_reg[28][25] , \partial_reg[28][24] , \partial_reg[28][23] , \partial_reg[28][22] , 
    \partial_reg[28][21] , \partial_reg[28][20] , \partial_reg[28][19] , \partial_reg[28][18] , 
    \partial_reg[28][17] , \partial_reg[28][16] , \partial_reg[28][15] , \partial_reg[28][14] , 
    \partial_reg[28][13] , \partial_reg[28][12] , \partial_reg[28][11] , \partial_reg[28][10] , 
    \partial_reg[28][9] , \partial_reg[28][8] , \partial_reg[28][7] , \partial_reg[28][6] , 
    \partial_reg[28][5] , \partial_reg[28][4] , \partial_reg[28][3] , \partial_reg[28][2] , 
    \partial_reg[28][1] , \partial_reg[28][0] }));
PartialAdder__1_2514 genblk1_25_p2 (.c1 ({\c1[25][31] , \c1[25][30] , \c1[25][29] , 
    \c1[25][28] , \c1[25][27] , \c1[25][26] , \c1[25][25] , \c1[25][24] , \c1[25][23] , 
    \c1[25][22] , \c1[25][21] , \c1[25][20] , \c1[25][19] , \c1[25][18] , \c1[25][17] , 
    \c1[25][16] , \c1[25][15] , \c1[25][14] , \c1[25][13] , \c1[25][12] , \c1[25][11] , 
    \c1[25][10] , \c1[25][9] , \c1[25][8] , \c1[25][7] , \c1[25][6] , \c1[25][5] , 
    \c1[25][4] , \c1[25][3] , \c1[25][2] , \c1[25][1] , \c1[25][0] }), .s1 ({uc_74, 
    n_39_798, n_39_797, n_39_796, n_39_795, n_39_794, n_39_793, n_39_792, n_39_791, 
    n_39_790, n_39_789, n_39_788, n_39_787, n_39_786, n_39_785, n_39_784, n_39_783, 
    n_39_782, n_39_781, n_39_780, n_39_779, n_39_778, n_39_777, n_39_776, n_39_775, 
    n_39_774, n_39_773, n_39_772, n_39_771, n_39_770, n_39_769, n_39_768, n_24}), .a ({
    \partial_reg[26][31] , n_39_766, n_39_765, n_39_764, n_39_763, n_39_762, n_39_761, 
    n_39_760, n_39_759, n_39_758, n_39_757, n_39_756, n_39_755, n_39_754, n_39_753, 
    n_39_752, n_39_751, n_39_750, n_39_749, n_39_748, n_39_747, n_39_746, n_39_745, 
    n_39_744, n_39_743, n_39_742, n_39_741, n_39_740, n_39_739, n_39_738, n_39_737, 
    n_39_736, uc_72}), .b ({\c1[24][31] , \c1[24][30] , \c1[24][29] , \c1[24][28] , 
    \c1[24][27] , \c1[24][26] , \c1[24][25] , \c1[24][24] , \c1[24][23] , \c1[24][22] , 
    \c1[24][21] , \c1[24][20] , \c1[24][19] , \c1[24][18] , \c1[24][17] , \c1[24][16] , 
    \c1[24][15] , \c1[24][14] , \c1[24][13] , \c1[24][12] , \c1[24][11] , \c1[24][10] , 
    \c1[24][9] , \c1[24][8] , \c1[24][7] , \c1[24][6] , \c1[24][5] , \c1[24][4] , 
    \c1[24][3] , \c1[24][2] , \c1[24][1] , \c1[24][0] }), .c ({uc_73, \partial_reg[27][30] , 
    \partial_reg[27][29] , \partial_reg[27][28] , \partial_reg[27][27] , \partial_reg[27][26] , 
    \partial_reg[27][25] , \partial_reg[27][24] , \partial_reg[27][23] , \partial_reg[27][22] , 
    \partial_reg[27][21] , \partial_reg[27][20] , \partial_reg[27][19] , \partial_reg[27][18] , 
    \partial_reg[27][17] , \partial_reg[27][16] , \partial_reg[27][15] , \partial_reg[27][14] , 
    \partial_reg[27][13] , \partial_reg[27][12] , \partial_reg[27][11] , \partial_reg[27][10] , 
    \partial_reg[27][9] , \partial_reg[27][8] , \partial_reg[27][7] , \partial_reg[27][6] , 
    \partial_reg[27][5] , \partial_reg[27][4] , \partial_reg[27][3] , \partial_reg[27][2] , 
    \partial_reg[27][1] , \partial_reg[27][0] }));
PartialAdder__1_2417 genblk1_24_p2 (.c1 ({\c1[24][31] , \c1[24][30] , \c1[24][29] , 
    \c1[24][28] , \c1[24][27] , \c1[24][26] , \c1[24][25] , \c1[24][24] , \c1[24][23] , 
    \c1[24][22] , \c1[24][21] , \c1[24][20] , \c1[24][19] , \c1[24][18] , \c1[24][17] , 
    \c1[24][16] , \c1[24][15] , \c1[24][14] , \c1[24][13] , \c1[24][12] , \c1[24][11] , 
    \c1[24][10] , \c1[24][9] , \c1[24][8] , \c1[24][7] , \c1[24][6] , \c1[24][5] , 
    \c1[24][4] , \c1[24][3] , \c1[24][2] , \c1[24][1] , \c1[24][0] }), .s1 ({uc_71, 
    n_39_766, n_39_765, n_39_764, n_39_763, n_39_762, n_39_761, n_39_760, n_39_759, 
    n_39_758, n_39_757, n_39_756, n_39_755, n_39_754, n_39_753, n_39_752, n_39_751, 
    n_39_750, n_39_749, n_39_748, n_39_747, n_39_746, n_39_745, n_39_744, n_39_743, 
    n_39_742, n_39_741, n_39_740, n_39_739, n_39_738, n_39_737, n_39_736, n_23}), .a ({
    \partial_reg[25][31] , n_39_734, n_39_733, n_39_732, n_39_731, n_39_730, n_39_729, 
    n_39_728, n_39_727, n_39_726, n_39_725, n_39_724, n_39_723, n_39_722, n_39_721, 
    n_39_720, n_39_719, n_39_718, n_39_717, n_39_716, n_39_715, n_39_714, n_39_713, 
    n_39_712, n_39_711, n_39_710, n_39_709, n_39_708, n_39_707, n_39_706, n_39_705, 
    n_39_704, uc_69}), .b ({\c1[23][31] , \c1[23][30] , \c1[23][29] , \c1[23][28] , 
    \c1[23][27] , \c1[23][26] , \c1[23][25] , \c1[23][24] , \c1[23][23] , \c1[23][22] , 
    \c1[23][21] , \c1[23][20] , \c1[23][19] , \c1[23][18] , \c1[23][17] , \c1[23][16] , 
    \c1[23][15] , \c1[23][14] , \c1[23][13] , \c1[23][12] , \c1[23][11] , \c1[23][10] , 
    \c1[23][9] , \c1[23][8] , \c1[23][7] , \c1[23][6] , \c1[23][5] , \c1[23][4] , 
    \c1[23][3] , \c1[23][2] , \c1[23][1] , \c1[23][0] }), .c ({uc_70, \partial_reg[26][30] , 
    \partial_reg[26][29] , \partial_reg[26][28] , \partial_reg[26][27] , \partial_reg[26][26] , 
    \partial_reg[26][25] , \partial_reg[26][24] , \partial_reg[26][23] , \partial_reg[26][22] , 
    \partial_reg[26][21] , \partial_reg[26][20] , \partial_reg[26][19] , \partial_reg[26][18] , 
    \partial_reg[26][17] , \partial_reg[26][16] , \partial_reg[26][15] , \partial_reg[26][14] , 
    \partial_reg[26][13] , \partial_reg[26][12] , \partial_reg[26][11] , \partial_reg[26][10] , 
    \partial_reg[26][9] , \partial_reg[26][8] , \partial_reg[26][7] , \partial_reg[26][6] , 
    \partial_reg[26][5] , \partial_reg[26][4] , \partial_reg[26][3] , \partial_reg[26][2] , 
    \partial_reg[26][1] , \partial_reg[26][0] }));
PartialAdder__1_2320 genblk1_23_p2 (.c1 ({\c1[23][31] , \c1[23][30] , \c1[23][29] , 
    \c1[23][28] , \c1[23][27] , \c1[23][26] , \c1[23][25] , \c1[23][24] , \c1[23][23] , 
    \c1[23][22] , \c1[23][21] , \c1[23][20] , \c1[23][19] , \c1[23][18] , \c1[23][17] , 
    \c1[23][16] , \c1[23][15] , \c1[23][14] , \c1[23][13] , \c1[23][12] , \c1[23][11] , 
    \c1[23][10] , \c1[23][9] , \c1[23][8] , \c1[23][7] , \c1[23][6] , \c1[23][5] , 
    \c1[23][4] , \c1[23][3] , \c1[23][2] , \c1[23][1] , \c1[23][0] }), .s1 ({uc_68, 
    n_39_734, n_39_733, n_39_732, n_39_731, n_39_730, n_39_729, n_39_728, n_39_727, 
    n_39_726, n_39_725, n_39_724, n_39_723, n_39_722, n_39_721, n_39_720, n_39_719, 
    n_39_718, n_39_717, n_39_716, n_39_715, n_39_714, n_39_713, n_39_712, n_39_711, 
    n_39_710, n_39_709, n_39_708, n_39_707, n_39_706, n_39_705, n_39_704, n_22}), .a ({
    \partial_reg[24][31] , n_39_702, n_39_701, n_39_700, n_39_699, n_39_698, n_39_697, 
    n_39_696, n_39_695, n_39_694, n_39_693, n_39_692, n_39_691, n_39_690, n_39_689, 
    n_39_688, n_39_687, n_39_686, n_39_685, n_39_684, n_39_683, n_39_682, n_39_681, 
    n_39_680, n_39_679, n_39_678, n_39_677, n_39_676, n_39_675, n_39_674, n_39_673, 
    n_39_672, uc_66}), .b ({\c1[22][31] , \c1[22][30] , \c1[22][29] , \c1[22][28] , 
    \c1[22][27] , \c1[22][26] , \c1[22][25] , \c1[22][24] , \c1[22][23] , \c1[22][22] , 
    \c1[22][21] , \c1[22][20] , \c1[22][19] , \c1[22][18] , \c1[22][17] , \c1[22][16] , 
    \c1[22][15] , \c1[22][14] , \c1[22][13] , \c1[22][12] , \c1[22][11] , \c1[22][10] , 
    \c1[22][9] , \c1[22][8] , \c1[22][7] , \c1[22][6] , \c1[22][5] , \c1[22][4] , 
    \c1[22][3] , \c1[22][2] , \c1[22][1] , \c1[22][0] }), .c ({uc_67, \partial_reg[25][30] , 
    \partial_reg[25][29] , \partial_reg[25][28] , \partial_reg[25][27] , \partial_reg[25][26] , 
    \partial_reg[25][25] , \partial_reg[25][24] , \partial_reg[25][23] , \partial_reg[25][22] , 
    \partial_reg[25][21] , \partial_reg[25][20] , \partial_reg[25][19] , \partial_reg[25][18] , 
    \partial_reg[25][17] , \partial_reg[25][16] , \partial_reg[25][15] , \partial_reg[25][14] , 
    \partial_reg[25][13] , \partial_reg[25][12] , \partial_reg[25][11] , \partial_reg[25][10] , 
    \partial_reg[25][9] , \partial_reg[25][8] , \partial_reg[25][7] , \partial_reg[25][6] , 
    \partial_reg[25][5] , \partial_reg[25][4] , \partial_reg[25][3] , \partial_reg[25][2] , 
    \partial_reg[25][1] , \partial_reg[25][0] }));
PartialAdder__1_2223 genblk1_22_p2 (.c1 ({\c1[22][31] , \c1[22][30] , \c1[22][29] , 
    \c1[22][28] , \c1[22][27] , \c1[22][26] , \c1[22][25] , \c1[22][24] , \c1[22][23] , 
    \c1[22][22] , \c1[22][21] , \c1[22][20] , \c1[22][19] , \c1[22][18] , \c1[22][17] , 
    \c1[22][16] , \c1[22][15] , \c1[22][14] , \c1[22][13] , \c1[22][12] , \c1[22][11] , 
    \c1[22][10] , \c1[22][9] , \c1[22][8] , \c1[22][7] , \c1[22][6] , \c1[22][5] , 
    \c1[22][4] , \c1[22][3] , \c1[22][2] , \c1[22][1] , \c1[22][0] }), .s1 ({uc_65, 
    n_39_702, n_39_701, n_39_700, n_39_699, n_39_698, n_39_697, n_39_696, n_39_695, 
    n_39_694, n_39_693, n_39_692, n_39_691, n_39_690, n_39_689, n_39_688, n_39_687, 
    n_39_686, n_39_685, n_39_684, n_39_683, n_39_682, n_39_681, n_39_680, n_39_679, 
    n_39_678, n_39_677, n_39_676, n_39_675, n_39_674, n_39_673, n_39_672, n_21}), .a ({
    \partial_reg[23][31] , n_39_670, n_39_669, n_39_668, n_39_667, n_39_666, n_39_665, 
    n_39_664, n_39_663, n_39_662, n_39_661, n_39_660, n_39_659, n_39_658, n_39_657, 
    n_39_656, n_39_655, n_39_654, n_39_653, n_39_652, n_39_651, n_39_650, n_39_649, 
    n_39_648, n_39_647, n_39_646, n_39_645, n_39_644, n_39_643, n_39_642, n_39_641, 
    n_39_640, uc_63}), .b ({\c1[21][31] , \c1[21][30] , \c1[21][29] , \c1[21][28] , 
    \c1[21][27] , \c1[21][26] , \c1[21][25] , \c1[21][24] , \c1[21][23] , \c1[21][22] , 
    \c1[21][21] , \c1[21][20] , \c1[21][19] , \c1[21][18] , \c1[21][17] , \c1[21][16] , 
    \c1[21][15] , \c1[21][14] , \c1[21][13] , \c1[21][12] , \c1[21][11] , \c1[21][10] , 
    \c1[21][9] , \c1[21][8] , \c1[21][7] , \c1[21][6] , \c1[21][5] , \c1[21][4] , 
    \c1[21][3] , \c1[21][2] , \c1[21][1] , \c1[21][0] }), .c ({uc_64, \partial_reg[24][30] , 
    \partial_reg[24][29] , \partial_reg[24][28] , \partial_reg[24][27] , \partial_reg[24][26] , 
    \partial_reg[24][25] , \partial_reg[24][24] , \partial_reg[24][23] , \partial_reg[24][22] , 
    \partial_reg[24][21] , \partial_reg[24][20] , \partial_reg[24][19] , \partial_reg[24][18] , 
    \partial_reg[24][17] , \partial_reg[24][16] , \partial_reg[24][15] , \partial_reg[24][14] , 
    \partial_reg[24][13] , \partial_reg[24][12] , \partial_reg[24][11] , \partial_reg[24][10] , 
    \partial_reg[24][9] , \partial_reg[24][8] , \partial_reg[24][7] , \partial_reg[24][6] , 
    \partial_reg[24][5] , \partial_reg[24][4] , \partial_reg[24][3] , \partial_reg[24][2] , 
    \partial_reg[24][1] , \partial_reg[24][0] }));
PartialAdder__1_2126 genblk1_21_p2 (.c1 ({\c1[21][31] , \c1[21][30] , \c1[21][29] , 
    \c1[21][28] , \c1[21][27] , \c1[21][26] , \c1[21][25] , \c1[21][24] , \c1[21][23] , 
    \c1[21][22] , \c1[21][21] , \c1[21][20] , \c1[21][19] , \c1[21][18] , \c1[21][17] , 
    \c1[21][16] , \c1[21][15] , \c1[21][14] , \c1[21][13] , \c1[21][12] , \c1[21][11] , 
    \c1[21][10] , \c1[21][9] , \c1[21][8] , \c1[21][7] , \c1[21][6] , \c1[21][5] , 
    \c1[21][4] , \c1[21][3] , \c1[21][2] , \c1[21][1] , \c1[21][0] }), .s1 ({uc_62, 
    n_39_670, n_39_669, n_39_668, n_39_667, n_39_666, n_39_665, n_39_664, n_39_663, 
    n_39_662, n_39_661, n_39_660, n_39_659, n_39_658, n_39_657, n_39_656, n_39_655, 
    n_39_654, n_39_653, n_39_652, n_39_651, n_39_650, n_39_649, n_39_648, n_39_647, 
    n_39_646, n_39_645, n_39_644, n_39_643, n_39_642, n_39_641, n_39_640, n_20}), .a ({
    \partial_reg[22][31] , n_39_638, n_39_637, n_39_636, n_39_635, n_39_634, n_39_633, 
    n_39_632, n_39_631, n_39_630, n_39_629, n_39_628, n_39_627, n_39_626, n_39_625, 
    n_39_624, n_39_623, n_39_622, n_39_621, n_39_620, n_39_619, n_39_618, n_39_617, 
    n_39_616, n_39_615, n_39_614, n_39_613, n_39_612, n_39_611, n_39_610, n_39_609, 
    n_39_608, uc_60}), .b ({\c1[20][31] , \c1[20][30] , \c1[20][29] , \c1[20][28] , 
    \c1[20][27] , \c1[20][26] , \c1[20][25] , \c1[20][24] , \c1[20][23] , \c1[20][22] , 
    \c1[20][21] , \c1[20][20] , \c1[20][19] , \c1[20][18] , \c1[20][17] , \c1[20][16] , 
    \c1[20][15] , \c1[20][14] , \c1[20][13] , \c1[20][12] , \c1[20][11] , \c1[20][10] , 
    \c1[20][9] , \c1[20][8] , \c1[20][7] , \c1[20][6] , \c1[20][5] , \c1[20][4] , 
    \c1[20][3] , \c1[20][2] , \c1[20][1] , \c1[20][0] }), .c ({uc_61, \partial_reg[23][30] , 
    \partial_reg[23][29] , \partial_reg[23][28] , \partial_reg[23][27] , \partial_reg[23][26] , 
    \partial_reg[23][25] , \partial_reg[23][24] , \partial_reg[23][23] , \partial_reg[23][22] , 
    \partial_reg[23][21] , \partial_reg[23][20] , \partial_reg[23][19] , \partial_reg[23][18] , 
    \partial_reg[23][17] , \partial_reg[23][16] , \partial_reg[23][15] , \partial_reg[23][14] , 
    \partial_reg[23][13] , \partial_reg[23][12] , \partial_reg[23][11] , \partial_reg[23][10] , 
    \partial_reg[23][9] , \partial_reg[23][8] , \partial_reg[23][7] , \partial_reg[23][6] , 
    \partial_reg[23][5] , \partial_reg[23][4] , \partial_reg[23][3] , \partial_reg[23][2] , 
    \partial_reg[23][1] , \partial_reg[23][0] }));
PartialAdder__1_2029 genblk1_20_p2 (.c1 ({\c1[20][31] , \c1[20][30] , \c1[20][29] , 
    \c1[20][28] , \c1[20][27] , \c1[20][26] , \c1[20][25] , \c1[20][24] , \c1[20][23] , 
    \c1[20][22] , \c1[20][21] , \c1[20][20] , \c1[20][19] , \c1[20][18] , \c1[20][17] , 
    \c1[20][16] , \c1[20][15] , \c1[20][14] , \c1[20][13] , \c1[20][12] , \c1[20][11] , 
    \c1[20][10] , \c1[20][9] , \c1[20][8] , \c1[20][7] , \c1[20][6] , \c1[20][5] , 
    \c1[20][4] , \c1[20][3] , \c1[20][2] , \c1[20][1] , \c1[20][0] }), .s1 ({uc_59, 
    n_39_638, n_39_637, n_39_636, n_39_635, n_39_634, n_39_633, n_39_632, n_39_631, 
    n_39_630, n_39_629, n_39_628, n_39_627, n_39_626, n_39_625, n_39_624, n_39_623, 
    n_39_622, n_39_621, n_39_620, n_39_619, n_39_618, n_39_617, n_39_616, n_39_615, 
    n_39_614, n_39_613, n_39_612, n_39_611, n_39_610, n_39_609, n_39_608, n_19}), .a ({
    \partial_reg[21][31] , n_39_606, n_39_605, n_39_604, n_39_603, n_39_602, n_39_601, 
    n_39_600, n_39_599, n_39_598, n_39_597, n_39_596, n_39_595, n_39_594, n_39_593, 
    n_39_592, n_39_591, n_39_590, n_39_589, n_39_588, n_39_587, n_39_586, n_39_585, 
    n_39_584, n_39_583, n_39_582, n_39_581, n_39_580, n_39_579, n_39_578, n_39_577, 
    n_39_576, uc_57}), .b ({\c1[19][31] , \c1[19][30] , \c1[19][29] , \c1[19][28] , 
    \c1[19][27] , \c1[19][26] , \c1[19][25] , \c1[19][24] , \c1[19][23] , \c1[19][22] , 
    \c1[19][21] , \c1[19][20] , \c1[19][19] , \c1[19][18] , \c1[19][17] , \c1[19][16] , 
    \c1[19][15] , \c1[19][14] , \c1[19][13] , \c1[19][12] , \c1[19][11] , \c1[19][10] , 
    \c1[19][9] , \c1[19][8] , \c1[19][7] , \c1[19][6] , \c1[19][5] , \c1[19][4] , 
    \c1[19][3] , \c1[19][2] , \c1[19][1] , \c1[19][0] }), .c ({uc_58, \partial_reg[22][30] , 
    \partial_reg[22][29] , \partial_reg[22][28] , \partial_reg[22][27] , \partial_reg[22][26] , 
    \partial_reg[22][25] , \partial_reg[22][24] , \partial_reg[22][23] , \partial_reg[22][22] , 
    \partial_reg[22][21] , \partial_reg[22][20] , \partial_reg[22][19] , \partial_reg[22][18] , 
    \partial_reg[22][17] , \partial_reg[22][16] , \partial_reg[22][15] , \partial_reg[22][14] , 
    \partial_reg[22][13] , \partial_reg[22][12] , \partial_reg[22][11] , \partial_reg[22][10] , 
    \partial_reg[22][9] , \partial_reg[22][8] , \partial_reg[22][7] , \partial_reg[22][6] , 
    \partial_reg[22][5] , \partial_reg[22][4] , \partial_reg[22][3] , \partial_reg[22][2] , 
    \partial_reg[22][1] , \partial_reg[22][0] }));
PartialAdder__1_1932 genblk1_19_p2 (.c1 ({\c1[19][31] , \c1[19][30] , \c1[19][29] , 
    \c1[19][28] , \c1[19][27] , \c1[19][26] , \c1[19][25] , \c1[19][24] , \c1[19][23] , 
    \c1[19][22] , \c1[19][21] , \c1[19][20] , \c1[19][19] , \c1[19][18] , \c1[19][17] , 
    \c1[19][16] , \c1[19][15] , \c1[19][14] , \c1[19][13] , \c1[19][12] , \c1[19][11] , 
    \c1[19][10] , \c1[19][9] , \c1[19][8] , \c1[19][7] , \c1[19][6] , \c1[19][5] , 
    \c1[19][4] , \c1[19][3] , \c1[19][2] , \c1[19][1] , \c1[19][0] }), .s1 ({uc_56, 
    n_39_606, n_39_605, n_39_604, n_39_603, n_39_602, n_39_601, n_39_600, n_39_599, 
    n_39_598, n_39_597, n_39_596, n_39_595, n_39_594, n_39_593, n_39_592, n_39_591, 
    n_39_590, n_39_589, n_39_588, n_39_587, n_39_586, n_39_585, n_39_584, n_39_583, 
    n_39_582, n_39_581, n_39_580, n_39_579, n_39_578, n_39_577, n_39_576, n_18}), .a ({
    \partial_reg[20][31] , n_39_574, n_39_573, n_39_572, n_39_571, n_39_570, n_39_569, 
    n_39_568, n_39_567, n_39_566, n_39_565, n_39_564, n_39_563, n_39_562, n_39_561, 
    n_39_560, n_39_559, n_39_558, n_39_557, n_39_556, n_39_555, n_39_554, n_39_553, 
    n_39_552, n_39_551, n_39_550, n_39_549, n_39_548, n_39_547, n_39_546, n_39_545, 
    n_39_544, uc_54}), .b ({\c1[18][31] , \c1[18][30] , \c1[18][29] , \c1[18][28] , 
    \c1[18][27] , \c1[18][26] , \c1[18][25] , \c1[18][24] , \c1[18][23] , \c1[18][22] , 
    \c1[18][21] , \c1[18][20] , \c1[18][19] , \c1[18][18] , \c1[18][17] , \c1[18][16] , 
    \c1[18][15] , \c1[18][14] , \c1[18][13] , \c1[18][12] , \c1[18][11] , \c1[18][10] , 
    \c1[18][9] , \c1[18][8] , \c1[18][7] , \c1[18][6] , \c1[18][5] , \c1[18][4] , 
    \c1[18][3] , \c1[18][2] , \c1[18][1] , \c1[18][0] }), .c ({uc_55, \partial_reg[21][30] , 
    \partial_reg[21][29] , \partial_reg[21][28] , \partial_reg[21][27] , \partial_reg[21][26] , 
    \partial_reg[21][25] , \partial_reg[21][24] , \partial_reg[21][23] , \partial_reg[21][22] , 
    \partial_reg[21][21] , \partial_reg[21][20] , \partial_reg[21][19] , \partial_reg[21][18] , 
    \partial_reg[21][17] , \partial_reg[21][16] , \partial_reg[21][15] , \partial_reg[21][14] , 
    \partial_reg[21][13] , \partial_reg[21][12] , \partial_reg[21][11] , \partial_reg[21][10] , 
    \partial_reg[21][9] , \partial_reg[21][8] , \partial_reg[21][7] , \partial_reg[21][6] , 
    \partial_reg[21][5] , \partial_reg[21][4] , \partial_reg[21][3] , \partial_reg[21][2] , 
    \partial_reg[21][1] , \partial_reg[21][0] }));
PartialAdder__1_1835 genblk1_18_p2 (.c1 ({\c1[18][31] , \c1[18][30] , \c1[18][29] , 
    \c1[18][28] , \c1[18][27] , \c1[18][26] , \c1[18][25] , \c1[18][24] , \c1[18][23] , 
    \c1[18][22] , \c1[18][21] , \c1[18][20] , \c1[18][19] , \c1[18][18] , \c1[18][17] , 
    \c1[18][16] , \c1[18][15] , \c1[18][14] , \c1[18][13] , \c1[18][12] , \c1[18][11] , 
    \c1[18][10] , \c1[18][9] , \c1[18][8] , \c1[18][7] , \c1[18][6] , \c1[18][5] , 
    \c1[18][4] , \c1[18][3] , \c1[18][2] , \c1[18][1] , \c1[18][0] }), .s1 ({uc_53, 
    n_39_574, n_39_573, n_39_572, n_39_571, n_39_570, n_39_569, n_39_568, n_39_567, 
    n_39_566, n_39_565, n_39_564, n_39_563, n_39_562, n_39_561, n_39_560, n_39_559, 
    n_39_558, n_39_557, n_39_556, n_39_555, n_39_554, n_39_553, n_39_552, n_39_551, 
    n_39_550, n_39_549, n_39_548, n_39_547, n_39_546, n_39_545, n_39_544, n_17}), .a ({
    \partial_reg[19][31] , n_39_542, n_39_541, n_39_540, n_39_539, n_39_538, n_39_537, 
    n_39_536, n_39_535, n_39_534, n_39_533, n_39_532, n_39_531, n_39_530, n_39_529, 
    n_39_528, n_39_527, n_39_526, n_39_525, n_39_524, n_39_523, n_39_522, n_39_521, 
    n_39_520, n_39_519, n_39_518, n_39_517, n_39_516, n_39_515, n_39_514, n_39_513, 
    n_39_512, uc_51}), .b ({\c1[17][31] , \c1[17][30] , \c1[17][29] , \c1[17][28] , 
    \c1[17][27] , \c1[17][26] , \c1[17][25] , \c1[17][24] , \c1[17][23] , \c1[17][22] , 
    \c1[17][21] , \c1[17][20] , \c1[17][19] , \c1[17][18] , \c1[17][17] , \c1[17][16] , 
    \c1[17][15] , \c1[17][14] , \c1[17][13] , \c1[17][12] , \c1[17][11] , \c1[17][10] , 
    \c1[17][9] , \c1[17][8] , \c1[17][7] , \c1[17][6] , \c1[17][5] , \c1[17][4] , 
    \c1[17][3] , \c1[17][2] , \c1[17][1] , \c1[17][0] }), .c ({uc_52, \partial_reg[20][30] , 
    \partial_reg[20][29] , \partial_reg[20][28] , \partial_reg[20][27] , \partial_reg[20][26] , 
    \partial_reg[20][25] , \partial_reg[20][24] , \partial_reg[20][23] , \partial_reg[20][22] , 
    \partial_reg[20][21] , \partial_reg[20][20] , \partial_reg[20][19] , \partial_reg[20][18] , 
    \partial_reg[20][17] , \partial_reg[20][16] , \partial_reg[20][15] , \partial_reg[20][14] , 
    \partial_reg[20][13] , \partial_reg[20][12] , \partial_reg[20][11] , \partial_reg[20][10] , 
    \partial_reg[20][9] , \partial_reg[20][8] , \partial_reg[20][7] , \partial_reg[20][6] , 
    \partial_reg[20][5] , \partial_reg[20][4] , \partial_reg[20][3] , \partial_reg[20][2] , 
    \partial_reg[20][1] , \partial_reg[20][0] }));
PartialAdder__1_1738 genblk1_17_p2 (.c1 ({\c1[17][31] , \c1[17][30] , \c1[17][29] , 
    \c1[17][28] , \c1[17][27] , \c1[17][26] , \c1[17][25] , \c1[17][24] , \c1[17][23] , 
    \c1[17][22] , \c1[17][21] , \c1[17][20] , \c1[17][19] , \c1[17][18] , \c1[17][17] , 
    \c1[17][16] , \c1[17][15] , \c1[17][14] , \c1[17][13] , \c1[17][12] , \c1[17][11] , 
    \c1[17][10] , \c1[17][9] , \c1[17][8] , \c1[17][7] , \c1[17][6] , \c1[17][5] , 
    \c1[17][4] , \c1[17][3] , \c1[17][2] , \c1[17][1] , \c1[17][0] }), .s1 ({uc_50, 
    n_39_542, n_39_541, n_39_540, n_39_539, n_39_538, n_39_537, n_39_536, n_39_535, 
    n_39_534, n_39_533, n_39_532, n_39_531, n_39_530, n_39_529, n_39_528, n_39_527, 
    n_39_526, n_39_525, n_39_524, n_39_523, n_39_522, n_39_521, n_39_520, n_39_519, 
    n_39_518, n_39_517, n_39_516, n_39_515, n_39_514, n_39_513, n_39_512, n_16}), .a ({
    \partial_reg[18][31] , n_39_510, n_39_509, n_39_508, n_39_507, n_39_506, n_39_505, 
    n_39_504, n_39_503, n_39_502, n_39_501, n_39_500, n_39_499, n_39_498, n_39_497, 
    n_39_496, n_39_495, n_39_494, n_39_493, n_39_492, n_39_491, n_39_490, n_39_489, 
    n_39_488, n_39_487, n_39_486, n_39_485, n_39_484, n_39_483, n_39_482, n_39_481, 
    n_39_480, uc_48}), .b ({\c1[16][31] , \c1[16][30] , \c1[16][29] , \c1[16][28] , 
    \c1[16][27] , \c1[16][26] , \c1[16][25] , \c1[16][24] , \c1[16][23] , \c1[16][22] , 
    \c1[16][21] , \c1[16][20] , \c1[16][19] , \c1[16][18] , \c1[16][17] , \c1[16][16] , 
    \c1[16][15] , \c1[16][14] , \c1[16][13] , \c1[16][12] , \c1[16][11] , \c1[16][10] , 
    \c1[16][9] , \c1[16][8] , \c1[16][7] , \c1[16][6] , \c1[16][5] , \c1[16][4] , 
    \c1[16][3] , \c1[16][2] , \c1[16][1] , \c1[16][0] }), .c ({uc_49, \partial_reg[19][30] , 
    \partial_reg[19][29] , \partial_reg[19][28] , \partial_reg[19][27] , \partial_reg[19][26] , 
    \partial_reg[19][25] , \partial_reg[19][24] , \partial_reg[19][23] , \partial_reg[19][22] , 
    \partial_reg[19][21] , \partial_reg[19][20] , \partial_reg[19][19] , \partial_reg[19][18] , 
    \partial_reg[19][17] , \partial_reg[19][16] , \partial_reg[19][15] , \partial_reg[19][14] , 
    \partial_reg[19][13] , \partial_reg[19][12] , \partial_reg[19][11] , \partial_reg[19][10] , 
    \partial_reg[19][9] , \partial_reg[19][8] , \partial_reg[19][7] , \partial_reg[19][6] , 
    \partial_reg[19][5] , \partial_reg[19][4] , \partial_reg[19][3] , \partial_reg[19][2] , 
    \partial_reg[19][1] , \partial_reg[19][0] }));
PartialAdder__1_1641 genblk1_16_p2 (.c1 ({\c1[16][31] , \c1[16][30] , \c1[16][29] , 
    \c1[16][28] , \c1[16][27] , \c1[16][26] , \c1[16][25] , \c1[16][24] , \c1[16][23] , 
    \c1[16][22] , \c1[16][21] , \c1[16][20] , \c1[16][19] , \c1[16][18] , \c1[16][17] , 
    \c1[16][16] , \c1[16][15] , \c1[16][14] , \c1[16][13] , \c1[16][12] , \c1[16][11] , 
    \c1[16][10] , \c1[16][9] , \c1[16][8] , \c1[16][7] , \c1[16][6] , \c1[16][5] , 
    \c1[16][4] , \c1[16][3] , \c1[16][2] , \c1[16][1] , \c1[16][0] }), .s1 ({uc_47, 
    n_39_510, n_39_509, n_39_508, n_39_507, n_39_506, n_39_505, n_39_504, n_39_503, 
    n_39_502, n_39_501, n_39_500, n_39_499, n_39_498, n_39_497, n_39_496, n_39_495, 
    n_39_494, n_39_493, n_39_492, n_39_491, n_39_490, n_39_489, n_39_488, n_39_487, 
    n_39_486, n_39_485, n_39_484, n_39_483, n_39_482, n_39_481, n_39_480, n_15}), .a ({
    \partial_reg[17][31] , n_39_478, n_39_477, n_39_476, n_39_475, n_39_474, n_39_473, 
    n_39_472, n_39_471, n_39_470, n_39_469, n_39_468, n_39_467, n_39_466, n_39_465, 
    n_39_464, n_39_463, n_39_462, n_39_461, n_39_460, n_39_459, n_39_458, n_39_457, 
    n_39_456, n_39_455, n_39_454, n_39_453, n_39_452, n_39_451, n_39_450, n_39_449, 
    n_39_448, uc_45}), .b ({\c1[15][31] , \c1[15][30] , \c1[15][29] , \c1[15][28] , 
    \c1[15][27] , \c1[15][26] , \c1[15][25] , \c1[15][24] , \c1[15][23] , \c1[15][22] , 
    \c1[15][21] , \c1[15][20] , \c1[15][19] , \c1[15][18] , \c1[15][17] , \c1[15][16] , 
    \c1[15][15] , \c1[15][14] , \c1[15][13] , \c1[15][12] , \c1[15][11] , \c1[15][10] , 
    \c1[15][9] , \c1[15][8] , \c1[15][7] , \c1[15][6] , \c1[15][5] , \c1[15][4] , 
    \c1[15][3] , \c1[15][2] , \c1[15][1] , \c1[15][0] }), .c ({uc_46, \partial_reg[18][30] , 
    \partial_reg[18][29] , \partial_reg[18][28] , \partial_reg[18][27] , \partial_reg[18][26] , 
    \partial_reg[18][25] , \partial_reg[18][24] , \partial_reg[18][23] , \partial_reg[18][22] , 
    \partial_reg[18][21] , \partial_reg[18][20] , \partial_reg[18][19] , \partial_reg[18][18] , 
    \partial_reg[18][17] , \partial_reg[18][16] , \partial_reg[18][15] , \partial_reg[18][14] , 
    \partial_reg[18][13] , \partial_reg[18][12] , \partial_reg[18][11] , \partial_reg[18][10] , 
    \partial_reg[18][9] , \partial_reg[18][8] , \partial_reg[18][7] , \partial_reg[18][6] , 
    \partial_reg[18][5] , \partial_reg[18][4] , \partial_reg[18][3] , \partial_reg[18][2] , 
    \partial_reg[18][1] , \partial_reg[18][0] }));
PartialAdder__1_1544 genblk1_15_p2 (.c1 ({\c1[15][31] , \c1[15][30] , \c1[15][29] , 
    \c1[15][28] , \c1[15][27] , \c1[15][26] , \c1[15][25] , \c1[15][24] , \c1[15][23] , 
    \c1[15][22] , \c1[15][21] , \c1[15][20] , \c1[15][19] , \c1[15][18] , \c1[15][17] , 
    \c1[15][16] , \c1[15][15] , \c1[15][14] , \c1[15][13] , \c1[15][12] , \c1[15][11] , 
    \c1[15][10] , \c1[15][9] , \c1[15][8] , \c1[15][7] , \c1[15][6] , \c1[15][5] , 
    \c1[15][4] , \c1[15][3] , \c1[15][2] , \c1[15][1] , \c1[15][0] }), .s1 ({uc_44, 
    n_39_478, n_39_477, n_39_476, n_39_475, n_39_474, n_39_473, n_39_472, n_39_471, 
    n_39_470, n_39_469, n_39_468, n_39_467, n_39_466, n_39_465, n_39_464, n_39_463, 
    n_39_462, n_39_461, n_39_460, n_39_459, n_39_458, n_39_457, n_39_456, n_39_455, 
    n_39_454, n_39_453, n_39_452, n_39_451, n_39_450, n_39_449, n_39_448, n_14}), .a ({
    \partial_reg[16][31] , n_39_446, n_39_445, n_39_444, n_39_443, n_39_442, n_39_441, 
    n_39_440, n_39_439, n_39_438, n_39_437, n_39_436, n_39_435, n_39_434, n_39_433, 
    n_39_432, n_39_431, n_39_430, n_39_429, n_39_428, n_39_427, n_39_426, n_39_425, 
    n_39_424, n_39_423, n_39_422, n_39_421, n_39_420, n_39_419, n_39_418, n_39_417, 
    n_39_416, uc_42}), .b ({\c1[14][31] , \c1[14][30] , \c1[14][29] , \c1[14][28] , 
    \c1[14][27] , \c1[14][26] , \c1[14][25] , \c1[14][24] , \c1[14][23] , \c1[14][22] , 
    \c1[14][21] , \c1[14][20] , \c1[14][19] , \c1[14][18] , \c1[14][17] , \c1[14][16] , 
    \c1[14][15] , \c1[14][14] , \c1[14][13] , \c1[14][12] , \c1[14][11] , \c1[14][10] , 
    \c1[14][9] , \c1[14][8] , \c1[14][7] , \c1[14][6] , \c1[14][5] , \c1[14][4] , 
    \c1[14][3] , \c1[14][2] , \c1[14][1] , \c1[14][0] }), .c ({uc_43, \partial_reg[17][30] , 
    \partial_reg[17][29] , \partial_reg[17][28] , \partial_reg[17][27] , \partial_reg[17][26] , 
    \partial_reg[17][25] , \partial_reg[17][24] , \partial_reg[17][23] , \partial_reg[17][22] , 
    \partial_reg[17][21] , \partial_reg[17][20] , \partial_reg[17][19] , \partial_reg[17][18] , 
    \partial_reg[17][17] , \partial_reg[17][16] , \partial_reg[17][15] , \partial_reg[17][14] , 
    \partial_reg[17][13] , \partial_reg[17][12] , \partial_reg[17][11] , \partial_reg[17][10] , 
    \partial_reg[17][9] , \partial_reg[17][8] , \partial_reg[17][7] , \partial_reg[17][6] , 
    \partial_reg[17][5] , \partial_reg[17][4] , \partial_reg[17][3] , \partial_reg[17][2] , 
    \partial_reg[17][1] , \partial_reg[17][0] }));
PartialAdder__1_1447 genblk1_14_p2 (.c1 ({\c1[14][31] , \c1[14][30] , \c1[14][29] , 
    \c1[14][28] , \c1[14][27] , \c1[14][26] , \c1[14][25] , \c1[14][24] , \c1[14][23] , 
    \c1[14][22] , \c1[14][21] , \c1[14][20] , \c1[14][19] , \c1[14][18] , \c1[14][17] , 
    \c1[14][16] , \c1[14][15] , \c1[14][14] , \c1[14][13] , \c1[14][12] , \c1[14][11] , 
    \c1[14][10] , \c1[14][9] , \c1[14][8] , \c1[14][7] , \c1[14][6] , \c1[14][5] , 
    \c1[14][4] , \c1[14][3] , \c1[14][2] , \c1[14][1] , \c1[14][0] }), .s1 ({uc_41, 
    n_39_446, n_39_445, n_39_444, n_39_443, n_39_442, n_39_441, n_39_440, n_39_439, 
    n_39_438, n_39_437, n_39_436, n_39_435, n_39_434, n_39_433, n_39_432, n_39_431, 
    n_39_430, n_39_429, n_39_428, n_39_427, n_39_426, n_39_425, n_39_424, n_39_423, 
    n_39_422, n_39_421, n_39_420, n_39_419, n_39_418, n_39_417, n_39_416, n_13}), .a ({
    \partial_reg[15][31] , n_39_414, n_39_413, n_39_412, n_39_411, n_39_410, n_39_409, 
    n_39_408, n_39_407, n_39_406, n_39_405, n_39_404, n_39_403, n_39_402, n_39_401, 
    n_39_400, n_39_399, n_39_398, n_39_397, n_39_396, n_39_395, n_39_394, n_39_393, 
    n_39_392, n_39_391, n_39_390, n_39_389, n_39_388, n_39_387, n_39_386, n_39_385, 
    n_39_384, uc_39}), .b ({\c1[13][31] , \c1[13][30] , \c1[13][29] , \c1[13][28] , 
    \c1[13][27] , \c1[13][26] , \c1[13][25] , \c1[13][24] , \c1[13][23] , \c1[13][22] , 
    \c1[13][21] , \c1[13][20] , \c1[13][19] , \c1[13][18] , \c1[13][17] , \c1[13][16] , 
    \c1[13][15] , \c1[13][14] , \c1[13][13] , \c1[13][12] , \c1[13][11] , \c1[13][10] , 
    \c1[13][9] , \c1[13][8] , \c1[13][7] , \c1[13][6] , \c1[13][5] , \c1[13][4] , 
    \c1[13][3] , \c1[13][2] , \c1[13][1] , \c1[13][0] }), .c ({uc_40, \partial_reg[16][30] , 
    \partial_reg[16][29] , \partial_reg[16][28] , \partial_reg[16][27] , \partial_reg[16][26] , 
    \partial_reg[16][25] , \partial_reg[16][24] , \partial_reg[16][23] , \partial_reg[16][22] , 
    \partial_reg[16][21] , \partial_reg[16][20] , \partial_reg[16][19] , \partial_reg[16][18] , 
    \partial_reg[16][17] , \partial_reg[16][16] , \partial_reg[16][15] , \partial_reg[16][14] , 
    \partial_reg[16][13] , \partial_reg[16][12] , \partial_reg[16][11] , \partial_reg[16][10] , 
    \partial_reg[16][9] , \partial_reg[16][8] , \partial_reg[16][7] , \partial_reg[16][6] , 
    \partial_reg[16][5] , \partial_reg[16][4] , \partial_reg[16][3] , \partial_reg[16][2] , 
    \partial_reg[16][1] , \partial_reg[16][0] }));
PartialAdder__1_1350 genblk1_13_p2 (.c1 ({\c1[13][31] , \c1[13][30] , \c1[13][29] , 
    \c1[13][28] , \c1[13][27] , \c1[13][26] , \c1[13][25] , \c1[13][24] , \c1[13][23] , 
    \c1[13][22] , \c1[13][21] , \c1[13][20] , \c1[13][19] , \c1[13][18] , \c1[13][17] , 
    \c1[13][16] , \c1[13][15] , \c1[13][14] , \c1[13][13] , \c1[13][12] , \c1[13][11] , 
    \c1[13][10] , \c1[13][9] , \c1[13][8] , \c1[13][7] , \c1[13][6] , \c1[13][5] , 
    \c1[13][4] , \c1[13][3] , \c1[13][2] , \c1[13][1] , \c1[13][0] }), .s1 ({uc_38, 
    n_39_414, n_39_413, n_39_412, n_39_411, n_39_410, n_39_409, n_39_408, n_39_407, 
    n_39_406, n_39_405, n_39_404, n_39_403, n_39_402, n_39_401, n_39_400, n_39_399, 
    n_39_398, n_39_397, n_39_396, n_39_395, n_39_394, n_39_393, n_39_392, n_39_391, 
    n_39_390, n_39_389, n_39_388, n_39_387, n_39_386, n_39_385, n_39_384, n_12}), .a ({
    \partial_reg[14][31] , n_39_382, n_39_381, n_39_380, n_39_379, n_39_378, n_39_377, 
    n_39_376, n_39_375, n_39_374, n_39_373, n_39_372, n_39_371, n_39_370, n_39_369, 
    n_39_368, n_39_367, n_39_366, n_39_365, n_39_364, n_39_363, n_39_362, n_39_361, 
    n_39_360, n_39_359, n_39_358, n_39_357, n_39_356, n_39_355, n_39_354, n_39_353, 
    n_39_352, uc_36}), .b ({\c1[12][31] , \c1[12][30] , \c1[12][29] , \c1[12][28] , 
    \c1[12][27] , \c1[12][26] , \c1[12][25] , \c1[12][24] , \c1[12][23] , \c1[12][22] , 
    \c1[12][21] , \c1[12][20] , \c1[12][19] , \c1[12][18] , \c1[12][17] , \c1[12][16] , 
    \c1[12][15] , \c1[12][14] , \c1[12][13] , \c1[12][12] , \c1[12][11] , \c1[12][10] , 
    \c1[12][9] , \c1[12][8] , \c1[12][7] , \c1[12][6] , \c1[12][5] , \c1[12][4] , 
    \c1[12][3] , \c1[12][2] , \c1[12][1] , \c1[12][0] }), .c ({uc_37, \partial_reg[15][30] , 
    \partial_reg[15][29] , \partial_reg[15][28] , \partial_reg[15][27] , \partial_reg[15][26] , 
    \partial_reg[15][25] , \partial_reg[15][24] , \partial_reg[15][23] , \partial_reg[15][22] , 
    \partial_reg[15][21] , \partial_reg[15][20] , \partial_reg[15][19] , \partial_reg[15][18] , 
    \partial_reg[15][17] , \partial_reg[15][16] , \partial_reg[15][15] , \partial_reg[15][14] , 
    \partial_reg[15][13] , \partial_reg[15][12] , \partial_reg[15][11] , \partial_reg[15][10] , 
    \partial_reg[15][9] , \partial_reg[15][8] , \partial_reg[15][7] , \partial_reg[15][6] , 
    \partial_reg[15][5] , \partial_reg[15][4] , \partial_reg[15][3] , \partial_reg[15][2] , 
    \partial_reg[15][1] , \partial_reg[15][0] }));
PartialAdder__1_1253 genblk1_12_p2 (.c1 ({\c1[12][31] , \c1[12][30] , \c1[12][29] , 
    \c1[12][28] , \c1[12][27] , \c1[12][26] , \c1[12][25] , \c1[12][24] , \c1[12][23] , 
    \c1[12][22] , \c1[12][21] , \c1[12][20] , \c1[12][19] , \c1[12][18] , \c1[12][17] , 
    \c1[12][16] , \c1[12][15] , \c1[12][14] , \c1[12][13] , \c1[12][12] , \c1[12][11] , 
    \c1[12][10] , \c1[12][9] , \c1[12][8] , \c1[12][7] , \c1[12][6] , \c1[12][5] , 
    \c1[12][4] , \c1[12][3] , \c1[12][2] , \c1[12][1] , \c1[12][0] }), .s1 ({uc_35, 
    n_39_382, n_39_381, n_39_380, n_39_379, n_39_378, n_39_377, n_39_376, n_39_375, 
    n_39_374, n_39_373, n_39_372, n_39_371, n_39_370, n_39_369, n_39_368, n_39_367, 
    n_39_366, n_39_365, n_39_364, n_39_363, n_39_362, n_39_361, n_39_360, n_39_359, 
    n_39_358, n_39_357, n_39_356, n_39_355, n_39_354, n_39_353, n_39_352, n_11}), .a ({
    \partial_reg[13][31] , n_39_350, n_39_349, n_39_348, n_39_347, n_39_346, n_39_345, 
    n_39_344, n_39_343, n_39_342, n_39_341, n_39_340, n_39_339, n_39_338, n_39_337, 
    n_39_336, n_39_335, n_39_334, n_39_333, n_39_332, n_39_331, n_39_330, n_39_329, 
    n_39_328, n_39_327, n_39_326, n_39_325, n_39_324, n_39_323, n_39_322, n_39_321, 
    n_39_320, uc_33}), .b ({\c1[11][31] , \c1[11][30] , \c1[11][29] , \c1[11][28] , 
    \c1[11][27] , \c1[11][26] , \c1[11][25] , \c1[11][24] , \c1[11][23] , \c1[11][22] , 
    \c1[11][21] , \c1[11][20] , \c1[11][19] , \c1[11][18] , \c1[11][17] , \c1[11][16] , 
    \c1[11][15] , \c1[11][14] , \c1[11][13] , \c1[11][12] , \c1[11][11] , \c1[11][10] , 
    \c1[11][9] , \c1[11][8] , \c1[11][7] , \c1[11][6] , \c1[11][5] , \c1[11][4] , 
    \c1[11][3] , \c1[11][2] , \c1[11][1] , \c1[11][0] }), .c ({uc_34, \partial_reg[14][30] , 
    \partial_reg[14][29] , \partial_reg[14][28] , \partial_reg[14][27] , \partial_reg[14][26] , 
    \partial_reg[14][25] , \partial_reg[14][24] , \partial_reg[14][23] , \partial_reg[14][22] , 
    \partial_reg[14][21] , \partial_reg[14][20] , \partial_reg[14][19] , \partial_reg[14][18] , 
    \partial_reg[14][17] , \partial_reg[14][16] , \partial_reg[14][15] , \partial_reg[14][14] , 
    \partial_reg[14][13] , \partial_reg[14][12] , \partial_reg[14][11] , \partial_reg[14][10] , 
    \partial_reg[14][9] , \partial_reg[14][8] , \partial_reg[14][7] , \partial_reg[14][6] , 
    \partial_reg[14][5] , \partial_reg[14][4] , \partial_reg[14][3] , \partial_reg[14][2] , 
    \partial_reg[14][1] , \partial_reg[14][0] }));
PartialAdder__1_1156 genblk1_11_p2 (.c1 ({\c1[11][31] , \c1[11][30] , \c1[11][29] , 
    \c1[11][28] , \c1[11][27] , \c1[11][26] , \c1[11][25] , \c1[11][24] , \c1[11][23] , 
    \c1[11][22] , \c1[11][21] , \c1[11][20] , \c1[11][19] , \c1[11][18] , \c1[11][17] , 
    \c1[11][16] , \c1[11][15] , \c1[11][14] , \c1[11][13] , \c1[11][12] , \c1[11][11] , 
    \c1[11][10] , \c1[11][9] , \c1[11][8] , \c1[11][7] , \c1[11][6] , \c1[11][5] , 
    \c1[11][4] , \c1[11][3] , \c1[11][2] , \c1[11][1] , \c1[11][0] }), .s1 ({uc_32, 
    n_39_350, n_39_349, n_39_348, n_39_347, n_39_346, n_39_345, n_39_344, n_39_343, 
    n_39_342, n_39_341, n_39_340, n_39_339, n_39_338, n_39_337, n_39_336, n_39_335, 
    n_39_334, n_39_333, n_39_332, n_39_331, n_39_330, n_39_329, n_39_328, n_39_327, 
    n_39_326, n_39_325, n_39_324, n_39_323, n_39_322, n_39_321, n_39_320, n_10}), .a ({
    \partial_reg[12][31] , n_39_318, n_39_317, n_39_316, n_39_315, n_39_314, n_39_313, 
    n_39_312, n_39_311, n_39_310, n_39_309, n_39_308, n_39_307, n_39_306, n_39_305, 
    n_39_304, n_39_303, n_39_302, n_39_301, n_39_300, n_39_299, n_39_298, n_39_297, 
    n_39_296, n_39_295, n_39_294, n_39_293, n_39_292, n_39_291, n_39_290, n_39_289, 
    n_39_288, uc_30}), .b ({\c1[10][31] , \c1[10][30] , \c1[10][29] , \c1[10][28] , 
    \c1[10][27] , \c1[10][26] , \c1[10][25] , \c1[10][24] , \c1[10][23] , \c1[10][22] , 
    \c1[10][21] , \c1[10][20] , \c1[10][19] , \c1[10][18] , \c1[10][17] , \c1[10][16] , 
    \c1[10][15] , \c1[10][14] , \c1[10][13] , \c1[10][12] , \c1[10][11] , \c1[10][10] , 
    \c1[10][9] , \c1[10][8] , \c1[10][7] , \c1[10][6] , \c1[10][5] , \c1[10][4] , 
    \c1[10][3] , \c1[10][2] , \c1[10][1] , \c1[10][0] }), .c ({uc_31, \partial_reg[13][30] , 
    \partial_reg[13][29] , \partial_reg[13][28] , \partial_reg[13][27] , \partial_reg[13][26] , 
    \partial_reg[13][25] , \partial_reg[13][24] , \partial_reg[13][23] , \partial_reg[13][22] , 
    \partial_reg[13][21] , \partial_reg[13][20] , \partial_reg[13][19] , \partial_reg[13][18] , 
    \partial_reg[13][17] , \partial_reg[13][16] , \partial_reg[13][15] , \partial_reg[13][14] , 
    \partial_reg[13][13] , \partial_reg[13][12] , \partial_reg[13][11] , \partial_reg[13][10] , 
    \partial_reg[13][9] , \partial_reg[13][8] , \partial_reg[13][7] , \partial_reg[13][6] , 
    \partial_reg[13][5] , \partial_reg[13][4] , \partial_reg[13][3] , \partial_reg[13][2] , 
    \partial_reg[13][1] , \partial_reg[13][0] }));
PartialAdder__1_1059 genblk1_10_p2 (.c1 ({\c1[10][31] , \c1[10][30] , \c1[10][29] , 
    \c1[10][28] , \c1[10][27] , \c1[10][26] , \c1[10][25] , \c1[10][24] , \c1[10][23] , 
    \c1[10][22] , \c1[10][21] , \c1[10][20] , \c1[10][19] , \c1[10][18] , \c1[10][17] , 
    \c1[10][16] , \c1[10][15] , \c1[10][14] , \c1[10][13] , \c1[10][12] , \c1[10][11] , 
    \c1[10][10] , \c1[10][9] , \c1[10][8] , \c1[10][7] , \c1[10][6] , \c1[10][5] , 
    \c1[10][4] , \c1[10][3] , \c1[10][2] , \c1[10][1] , \c1[10][0] }), .s1 ({uc_29, 
    n_39_318, n_39_317, n_39_316, n_39_315, n_39_314, n_39_313, n_39_312, n_39_311, 
    n_39_310, n_39_309, n_39_308, n_39_307, n_39_306, n_39_305, n_39_304, n_39_303, 
    n_39_302, n_39_301, n_39_300, n_39_299, n_39_298, n_39_297, n_39_296, n_39_295, 
    n_39_294, n_39_293, n_39_292, n_39_291, n_39_290, n_39_289, n_39_288, n_9}), .a ({
    \partial_reg[11][31] , n_39_286, n_39_285, n_39_284, n_39_283, n_39_282, n_39_281, 
    n_39_280, n_39_279, n_39_278, n_39_277, n_39_276, n_39_275, n_39_274, n_39_273, 
    n_39_272, n_39_271, n_39_270, n_39_269, n_39_268, n_39_267, n_39_266, n_39_265, 
    n_39_264, n_39_263, n_39_262, n_39_261, n_39_260, n_39_259, n_39_258, n_39_257, 
    n_39_256, uc_27}), .b ({\c1[9][31] , \c1[9][30] , \c1[9][29] , \c1[9][28] , \c1[9][27] , 
    \c1[9][26] , \c1[9][25] , \c1[9][24] , \c1[9][23] , \c1[9][22] , \c1[9][21] , 
    \c1[9][20] , \c1[9][19] , \c1[9][18] , \c1[9][17] , \c1[9][16] , \c1[9][15] , 
    \c1[9][14] , \c1[9][13] , \c1[9][12] , \c1[9][11] , \c1[9][10] , \c1[9][9] , 
    \c1[9][8] , \c1[9][7] , \c1[9][6] , \c1[9][5] , \c1[9][4] , \c1[9][3] , \c1[9][2] , 
    \c1[9][1] , \c1[9][0] }), .c ({uc_28, \partial_reg[12][30] , \partial_reg[12][29] , 
    \partial_reg[12][28] , \partial_reg[12][27] , \partial_reg[12][26] , \partial_reg[12][25] , 
    \partial_reg[12][24] , \partial_reg[12][23] , \partial_reg[12][22] , \partial_reg[12][21] , 
    \partial_reg[12][20] , \partial_reg[12][19] , \partial_reg[12][18] , \partial_reg[12][17] , 
    \partial_reg[12][16] , \partial_reg[12][15] , \partial_reg[12][14] , \partial_reg[12][13] , 
    \partial_reg[12][12] , \partial_reg[12][11] , \partial_reg[12][10] , \partial_reg[12][9] , 
    \partial_reg[12][8] , \partial_reg[12][7] , \partial_reg[12][6] , \partial_reg[12][5] , 
    \partial_reg[12][4] , \partial_reg[12][3] , \partial_reg[12][2] , \partial_reg[12][1] , 
    \partial_reg[12][0] }));
PartialAdder__1_962 genblk1_9_p2 (.c1 ({\c1[9][31] , \c1[9][30] , \c1[9][29] , \c1[9][28] , 
    \c1[9][27] , \c1[9][26] , \c1[9][25] , \c1[9][24] , \c1[9][23] , \c1[9][22] , 
    \c1[9][21] , \c1[9][20] , \c1[9][19] , \c1[9][18] , \c1[9][17] , \c1[9][16] , 
    \c1[9][15] , \c1[9][14] , \c1[9][13] , \c1[9][12] , \c1[9][11] , \c1[9][10] , 
    \c1[9][9] , \c1[9][8] , \c1[9][7] , \c1[9][6] , \c1[9][5] , \c1[9][4] , \c1[9][3] , 
    \c1[9][2] , \c1[9][1] , \c1[9][0] }), .s1 ({uc_26, n_39_286, n_39_285, n_39_284, 
    n_39_283, n_39_282, n_39_281, n_39_280, n_39_279, n_39_278, n_39_277, n_39_276, 
    n_39_275, n_39_274, n_39_273, n_39_272, n_39_271, n_39_270, n_39_269, n_39_268, 
    n_39_267, n_39_266, n_39_265, n_39_264, n_39_263, n_39_262, n_39_261, n_39_260, 
    n_39_259, n_39_258, n_39_257, n_39_256, n_8}), .a ({\partial_reg[10][31] , n_39_254, 
    n_39_253, n_39_252, n_39_251, n_39_250, n_39_249, n_39_248, n_39_247, n_39_246, 
    n_39_245, n_39_244, n_39_243, n_39_242, n_39_241, n_39_240, n_39_239, n_39_238, 
    n_39_237, n_39_236, n_39_235, n_39_234, n_39_233, n_39_232, n_39_231, n_39_230, 
    n_39_229, n_39_228, n_39_227, n_39_226, n_39_225, n_39_224, uc_24}), .b ({\c1[8][31] , 
    \c1[8][30] , \c1[8][29] , \c1[8][28] , \c1[8][27] , \c1[8][26] , \c1[8][25] , 
    \c1[8][24] , \c1[8][23] , \c1[8][22] , \c1[8][21] , \c1[8][20] , \c1[8][19] , 
    \c1[8][18] , \c1[8][17] , \c1[8][16] , \c1[8][15] , \c1[8][14] , \c1[8][13] , 
    \c1[8][12] , \c1[8][11] , \c1[8][10] , \c1[8][9] , \c1[8][8] , \c1[8][7] , \c1[8][6] , 
    \c1[8][5] , \c1[8][4] , \c1[8][3] , \c1[8][2] , \c1[8][1] , \c1[8][0] }), .c ({
    uc_25, \partial_reg[11][30] , \partial_reg[11][29] , \partial_reg[11][28] , \partial_reg[11][27] , 
    \partial_reg[11][26] , \partial_reg[11][25] , \partial_reg[11][24] , \partial_reg[11][23] , 
    \partial_reg[11][22] , \partial_reg[11][21] , \partial_reg[11][20] , \partial_reg[11][19] , 
    \partial_reg[11][18] , \partial_reg[11][17] , \partial_reg[11][16] , \partial_reg[11][15] , 
    \partial_reg[11][14] , \partial_reg[11][13] , \partial_reg[11][12] , \partial_reg[11][11] , 
    \partial_reg[11][10] , \partial_reg[11][9] , \partial_reg[11][8] , \partial_reg[11][7] , 
    \partial_reg[11][6] , \partial_reg[11][5] , \partial_reg[11][4] , \partial_reg[11][3] , 
    \partial_reg[11][2] , \partial_reg[11][1] , \partial_reg[11][0] }));
PartialAdder__1_865 genblk1_8_p2 (.c1 ({\c1[8][31] , \c1[8][30] , \c1[8][29] , \c1[8][28] , 
    \c1[8][27] , \c1[8][26] , \c1[8][25] , \c1[8][24] , \c1[8][23] , \c1[8][22] , 
    \c1[8][21] , \c1[8][20] , \c1[8][19] , \c1[8][18] , \c1[8][17] , \c1[8][16] , 
    \c1[8][15] , \c1[8][14] , \c1[8][13] , \c1[8][12] , \c1[8][11] , \c1[8][10] , 
    \c1[8][9] , \c1[8][8] , \c1[8][7] , \c1[8][6] , \c1[8][5] , \c1[8][4] , \c1[8][3] , 
    \c1[8][2] , \c1[8][1] , \c1[8][0] }), .s1 ({uc_23, n_39_254, n_39_253, n_39_252, 
    n_39_251, n_39_250, n_39_249, n_39_248, n_39_247, n_39_246, n_39_245, n_39_244, 
    n_39_243, n_39_242, n_39_241, n_39_240, n_39_239, n_39_238, n_39_237, n_39_236, 
    n_39_235, n_39_234, n_39_233, n_39_232, n_39_231, n_39_230, n_39_229, n_39_228, 
    n_39_227, n_39_226, n_39_225, n_39_224, n_7}), .a ({\partial_reg[9][31] , n_39_222, 
    n_39_221, n_39_220, n_39_219, n_39_218, n_39_217, n_39_216, n_39_215, n_39_214, 
    n_39_213, n_39_212, n_39_211, n_39_210, n_39_209, n_39_208, n_39_207, n_39_206, 
    n_39_205, n_39_204, n_39_203, n_39_202, n_39_201, n_39_200, n_39_199, n_39_198, 
    n_39_197, n_39_196, n_39_195, n_39_194, n_39_193, n_39_192, uc_21}), .b ({\c1[7][31] , 
    \c1[7][30] , \c1[7][29] , \c1[7][28] , \c1[7][27] , \c1[7][26] , \c1[7][25] , 
    \c1[7][24] , \c1[7][23] , \c1[7][22] , \c1[7][21] , \c1[7][20] , \c1[7][19] , 
    \c1[7][18] , \c1[7][17] , \c1[7][16] , \c1[7][15] , \c1[7][14] , \c1[7][13] , 
    \c1[7][12] , \c1[7][11] , \c1[7][10] , \c1[7][9] , \c1[7][8] , \c1[7][7] , \c1[7][6] , 
    \c1[7][5] , \c1[7][4] , \c1[7][3] , \c1[7][2] , \c1[7][1] , \c1[7][0] }), .c ({
    uc_22, \partial_reg[10][30] , \partial_reg[10][29] , \partial_reg[10][28] , \partial_reg[10][27] , 
    \partial_reg[10][26] , \partial_reg[10][25] , \partial_reg[10][24] , \partial_reg[10][23] , 
    \partial_reg[10][22] , \partial_reg[10][21] , \partial_reg[10][20] , \partial_reg[10][19] , 
    \partial_reg[10][18] , \partial_reg[10][17] , \partial_reg[10][16] , \partial_reg[10][15] , 
    \partial_reg[10][14] , \partial_reg[10][13] , \partial_reg[10][12] , \partial_reg[10][11] , 
    \partial_reg[10][10] , \partial_reg[10][9] , \partial_reg[10][8] , \partial_reg[10][7] , 
    \partial_reg[10][6] , \partial_reg[10][5] , \partial_reg[10][4] , \partial_reg[10][3] , 
    \partial_reg[10][2] , \partial_reg[10][1] , \partial_reg[10][0] }));
PartialAdder__1_768 genblk1_7_p2 (.c1 ({\c1[7][31] , \c1[7][30] , \c1[7][29] , \c1[7][28] , 
    \c1[7][27] , \c1[7][26] , \c1[7][25] , \c1[7][24] , \c1[7][23] , \c1[7][22] , 
    \c1[7][21] , \c1[7][20] , \c1[7][19] , \c1[7][18] , \c1[7][17] , \c1[7][16] , 
    \c1[7][15] , \c1[7][14] , \c1[7][13] , \c1[7][12] , \c1[7][11] , \c1[7][10] , 
    \c1[7][9] , \c1[7][8] , \c1[7][7] , \c1[7][6] , \c1[7][5] , \c1[7][4] , \c1[7][3] , 
    \c1[7][2] , \c1[7][1] , \c1[7][0] }), .s1 ({uc_20, n_39_222, n_39_221, n_39_220, 
    n_39_219, n_39_218, n_39_217, n_39_216, n_39_215, n_39_214, n_39_213, n_39_212, 
    n_39_211, n_39_210, n_39_209, n_39_208, n_39_207, n_39_206, n_39_205, n_39_204, 
    n_39_203, n_39_202, n_39_201, n_39_200, n_39_199, n_39_198, n_39_197, n_39_196, 
    n_39_195, n_39_194, n_39_193, n_39_192, n_6}), .a ({\partial_reg[8][31] , n_39_190, 
    n_39_189, n_39_188, n_39_187, n_39_186, n_39_185, n_39_184, n_39_183, n_39_182, 
    n_39_181, n_39_180, n_39_179, n_39_178, n_39_177, n_39_176, n_39_175, n_39_174, 
    n_39_173, n_39_172, n_39_171, n_39_170, n_39_169, n_39_168, n_39_167, n_39_166, 
    n_39_165, n_39_164, n_39_163, n_39_162, n_39_161, n_39_160, uc_18}), .b ({\c1[6][31] , 
    \c1[6][30] , \c1[6][29] , \c1[6][28] , \c1[6][27] , \c1[6][26] , \c1[6][25] , 
    \c1[6][24] , \c1[6][23] , \c1[6][22] , \c1[6][21] , \c1[6][20] , \c1[6][19] , 
    \c1[6][18] , \c1[6][17] , \c1[6][16] , \c1[6][15] , \c1[6][14] , \c1[6][13] , 
    \c1[6][12] , \c1[6][11] , \c1[6][10] , \c1[6][9] , \c1[6][8] , \c1[6][7] , \c1[6][6] , 
    \c1[6][5] , \c1[6][4] , \c1[6][3] , \c1[6][2] , \c1[6][1] , \c1[6][0] }), .c ({
    uc_19, \partial_reg[9][30] , \partial_reg[9][29] , \partial_reg[9][28] , \partial_reg[9][27] , 
    \partial_reg[9][26] , \partial_reg[9][25] , \partial_reg[9][24] , \partial_reg[9][23] , 
    \partial_reg[9][22] , \partial_reg[9][21] , \partial_reg[9][20] , \partial_reg[9][19] , 
    \partial_reg[9][18] , \partial_reg[9][17] , \partial_reg[9][16] , \partial_reg[9][15] , 
    \partial_reg[9][14] , \partial_reg[9][13] , \partial_reg[9][12] , \partial_reg[9][11] , 
    \partial_reg[9][10] , \partial_reg[9][9] , \partial_reg[9][8] , \partial_reg[9][7] , 
    \partial_reg[9][6] , \partial_reg[9][5] , \partial_reg[9][4] , \partial_reg[9][3] , 
    \partial_reg[9][2] , \partial_reg[9][1] , \partial_reg[9][0] }));
PartialAdder__1_671 genblk1_6_p2 (.c1 ({\c1[6][31] , \c1[6][30] , \c1[6][29] , \c1[6][28] , 
    \c1[6][27] , \c1[6][26] , \c1[6][25] , \c1[6][24] , \c1[6][23] , \c1[6][22] , 
    \c1[6][21] , \c1[6][20] , \c1[6][19] , \c1[6][18] , \c1[6][17] , \c1[6][16] , 
    \c1[6][15] , \c1[6][14] , \c1[6][13] , \c1[6][12] , \c1[6][11] , \c1[6][10] , 
    \c1[6][9] , \c1[6][8] , \c1[6][7] , \c1[6][6] , \c1[6][5] , \c1[6][4] , \c1[6][3] , 
    \c1[6][2] , \c1[6][1] , \c1[6][0] }), .s1 ({uc_17, n_39_190, n_39_189, n_39_188, 
    n_39_187, n_39_186, n_39_185, n_39_184, n_39_183, n_39_182, n_39_181, n_39_180, 
    n_39_179, n_39_178, n_39_177, n_39_176, n_39_175, n_39_174, n_39_173, n_39_172, 
    n_39_171, n_39_170, n_39_169, n_39_168, n_39_167, n_39_166, n_39_165, n_39_164, 
    n_39_163, n_39_162, n_39_161, n_39_160, n_5}), .a ({\partial_reg[7][31] , n_39_158, 
    n_39_157, n_39_156, n_39_155, n_39_154, n_39_153, n_39_152, n_39_151, n_39_150, 
    n_39_149, n_39_148, n_39_147, n_39_146, n_39_145, n_39_144, n_39_143, n_39_142, 
    n_39_141, n_39_140, n_39_139, n_39_138, n_39_137, n_39_136, n_39_135, n_39_134, 
    n_39_133, n_39_132, n_39_131, n_39_130, n_39_129, n_39_128, uc_15}), .b ({\c1[5][31] , 
    \c1[5][30] , \c1[5][29] , \c1[5][28] , \c1[5][27] , \c1[5][26] , \c1[5][25] , 
    \c1[5][24] , \c1[5][23] , \c1[5][22] , \c1[5][21] , \c1[5][20] , \c1[5][19] , 
    \c1[5][18] , \c1[5][17] , \c1[5][16] , \c1[5][15] , \c1[5][14] , \c1[5][13] , 
    \c1[5][12] , \c1[5][11] , \c1[5][10] , \c1[5][9] , \c1[5][8] , \c1[5][7] , \c1[5][6] , 
    \c1[5][5] , \c1[5][4] , \c1[5][3] , \c1[5][2] , \c1[5][1] , \c1[5][0] }), .c ({
    uc_16, \partial_reg[8][30] , \partial_reg[8][29] , \partial_reg[8][28] , \partial_reg[8][27] , 
    \partial_reg[8][26] , \partial_reg[8][25] , \partial_reg[8][24] , \partial_reg[8][23] , 
    \partial_reg[8][22] , \partial_reg[8][21] , \partial_reg[8][20] , \partial_reg[8][19] , 
    \partial_reg[8][18] , \partial_reg[8][17] , \partial_reg[8][16] , \partial_reg[8][15] , 
    \partial_reg[8][14] , \partial_reg[8][13] , \partial_reg[8][12] , \partial_reg[8][11] , 
    \partial_reg[8][10] , \partial_reg[8][9] , \partial_reg[8][8] , \partial_reg[8][7] , 
    \partial_reg[8][6] , \partial_reg[8][5] , \partial_reg[8][4] , \partial_reg[8][3] , 
    \partial_reg[8][2] , \partial_reg[8][1] , \partial_reg[8][0] }));
PartialAdder__1_574 genblk1_5_p2 (.c1 ({\c1[5][31] , \c1[5][30] , \c1[5][29] , \c1[5][28] , 
    \c1[5][27] , \c1[5][26] , \c1[5][25] , \c1[5][24] , \c1[5][23] , \c1[5][22] , 
    \c1[5][21] , \c1[5][20] , \c1[5][19] , \c1[5][18] , \c1[5][17] , \c1[5][16] , 
    \c1[5][15] , \c1[5][14] , \c1[5][13] , \c1[5][12] , \c1[5][11] , \c1[5][10] , 
    \c1[5][9] , \c1[5][8] , \c1[5][7] , \c1[5][6] , \c1[5][5] , \c1[5][4] , \c1[5][3] , 
    \c1[5][2] , \c1[5][1] , \c1[5][0] }), .s1 ({uc_14, n_39_158, n_39_157, n_39_156, 
    n_39_155, n_39_154, n_39_153, n_39_152, n_39_151, n_39_150, n_39_149, n_39_148, 
    n_39_147, n_39_146, n_39_145, n_39_144, n_39_143, n_39_142, n_39_141, n_39_140, 
    n_39_139, n_39_138, n_39_137, n_39_136, n_39_135, n_39_134, n_39_133, n_39_132, 
    n_39_131, n_39_130, n_39_129, n_39_128, n_4}), .a ({\partial_reg[6][31] , n_39_126, 
    n_39_125, n_39_124, n_39_123, n_39_122, n_39_121, n_39_120, n_39_119, n_39_118, 
    n_39_117, n_39_116, n_39_115, n_39_114, n_39_113, n_39_112, n_39_111, n_39_110, 
    n_39_109, n_39_108, n_39_107, n_39_106, n_39_105, n_39_104, n_39_103, n_39_102, 
    n_39_101, n_39_100, n_39_99, n_39_98, n_39_97, n_39_96, uc_12}), .b ({\c1[4][31] , 
    \c1[4][30] , \c1[4][29] , \c1[4][28] , \c1[4][27] , \c1[4][26] , \c1[4][25] , 
    \c1[4][24] , \c1[4][23] , \c1[4][22] , \c1[4][21] , \c1[4][20] , \c1[4][19] , 
    \c1[4][18] , \c1[4][17] , \c1[4][16] , \c1[4][15] , \c1[4][14] , \c1[4][13] , 
    \c1[4][12] , \c1[4][11] , \c1[4][10] , \c1[4][9] , \c1[4][8] , \c1[4][7] , \c1[4][6] , 
    \c1[4][5] , \c1[4][4] , \c1[4][3] , \c1[4][2] , \c1[4][1] , \c1[4][0] }), .c ({
    uc_13, \partial_reg[7][30] , \partial_reg[7][29] , \partial_reg[7][28] , \partial_reg[7][27] , 
    \partial_reg[7][26] , \partial_reg[7][25] , \partial_reg[7][24] , \partial_reg[7][23] , 
    \partial_reg[7][22] , \partial_reg[7][21] , \partial_reg[7][20] , \partial_reg[7][19] , 
    \partial_reg[7][18] , \partial_reg[7][17] , \partial_reg[7][16] , \partial_reg[7][15] , 
    \partial_reg[7][14] , \partial_reg[7][13] , \partial_reg[7][12] , \partial_reg[7][11] , 
    \partial_reg[7][10] , \partial_reg[7][9] , \partial_reg[7][8] , \partial_reg[7][7] , 
    \partial_reg[7][6] , \partial_reg[7][5] , \partial_reg[7][4] , \partial_reg[7][3] , 
    \partial_reg[7][2] , \partial_reg[7][1] , \partial_reg[7][0] }));
PartialAdder__1_477 genblk1_4_p2 (.c1 ({\c1[4][31] , \c1[4][30] , \c1[4][29] , \c1[4][28] , 
    \c1[4][27] , \c1[4][26] , \c1[4][25] , \c1[4][24] , \c1[4][23] , \c1[4][22] , 
    \c1[4][21] , \c1[4][20] , \c1[4][19] , \c1[4][18] , \c1[4][17] , \c1[4][16] , 
    \c1[4][15] , \c1[4][14] , \c1[4][13] , \c1[4][12] , \c1[4][11] , \c1[4][10] , 
    \c1[4][9] , \c1[4][8] , \c1[4][7] , \c1[4][6] , \c1[4][5] , \c1[4][4] , \c1[4][3] , 
    \c1[4][2] , \c1[4][1] , \c1[4][0] }), .s1 ({uc_11, n_39_126, n_39_125, n_39_124, 
    n_39_123, n_39_122, n_39_121, n_39_120, n_39_119, n_39_118, n_39_117, n_39_116, 
    n_39_115, n_39_114, n_39_113, n_39_112, n_39_111, n_39_110, n_39_109, n_39_108, 
    n_39_107, n_39_106, n_39_105, n_39_104, n_39_103, n_39_102, n_39_101, n_39_100, 
    n_39_99, n_39_98, n_39_97, n_39_96, n_3}), .a ({\partial_reg[5][31] , n_39_94, 
    n_39_93, n_39_92, n_39_91, n_39_90, n_39_89, n_39_88, n_39_87, n_39_86, n_39_85, 
    n_39_84, n_39_83, n_39_82, n_39_81, n_39_80, n_39_79, n_39_78, n_39_77, n_39_76, 
    n_39_75, n_39_74, n_39_73, n_39_72, n_39_71, n_39_70, n_39_69, n_39_68, n_39_67, 
    n_39_66, n_39_65, n_39_64, uc_9}), .b ({\c1[3][31] , \c1[3][30] , \c1[3][29] , 
    \c1[3][28] , \c1[3][27] , \c1[3][26] , \c1[3][25] , \c1[3][24] , \c1[3][23] , 
    \c1[3][22] , \c1[3][21] , \c1[3][20] , \c1[3][19] , \c1[3][18] , \c1[3][17] , 
    \c1[3][16] , \c1[3][15] , \c1[3][14] , \c1[3][13] , \c1[3][12] , \c1[3][11] , 
    \c1[3][10] , \c1[3][9] , \c1[3][8] , \c1[3][7] , \c1[3][6] , \c1[3][5] , \c1[3][4] , 
    \c1[3][3] , \c1[3][2] , \c1[3][1] , \c1[3][0] }), .c ({uc_10, \partial_reg[6][30] , 
    \partial_reg[6][29] , \partial_reg[6][28] , \partial_reg[6][27] , \partial_reg[6][26] , 
    \partial_reg[6][25] , \partial_reg[6][24] , \partial_reg[6][23] , \partial_reg[6][22] , 
    \partial_reg[6][21] , \partial_reg[6][20] , \partial_reg[6][19] , \partial_reg[6][18] , 
    \partial_reg[6][17] , \partial_reg[6][16] , \partial_reg[6][15] , \partial_reg[6][14] , 
    \partial_reg[6][13] , \partial_reg[6][12] , \partial_reg[6][11] , \partial_reg[6][10] , 
    \partial_reg[6][9] , \partial_reg[6][8] , \partial_reg[6][7] , \partial_reg[6][6] , 
    \partial_reg[6][5] , \partial_reg[6][4] , \partial_reg[6][3] , \partial_reg[6][2] , 
    \partial_reg[6][1] , \partial_reg[6][0] }));
PartialAdder__1_380 genblk1_3_p2 (.c1 ({\c1[3][31] , \c1[3][30] , \c1[3][29] , \c1[3][28] , 
    \c1[3][27] , \c1[3][26] , \c1[3][25] , \c1[3][24] , \c1[3][23] , \c1[3][22] , 
    \c1[3][21] , \c1[3][20] , \c1[3][19] , \c1[3][18] , \c1[3][17] , \c1[3][16] , 
    \c1[3][15] , \c1[3][14] , \c1[3][13] , \c1[3][12] , \c1[3][11] , \c1[3][10] , 
    \c1[3][9] , \c1[3][8] , \c1[3][7] , \c1[3][6] , \c1[3][5] , \c1[3][4] , \c1[3][3] , 
    \c1[3][2] , \c1[3][1] , \c1[3][0] }), .s1 ({uc_8, n_39_94, n_39_93, n_39_92, 
    n_39_91, n_39_90, n_39_89, n_39_88, n_39_87, n_39_86, n_39_85, n_39_84, n_39_83, 
    n_39_82, n_39_81, n_39_80, n_39_79, n_39_78, n_39_77, n_39_76, n_39_75, n_39_74, 
    n_39_73, n_39_72, n_39_71, n_39_70, n_39_69, n_39_68, n_39_67, n_39_66, n_39_65, 
    n_39_64, n_2}), .a ({\partial_reg[4][31] , n_39_62, n_39_61, n_39_60, n_39_59, 
    n_39_58, n_39_57, n_39_56, n_39_55, n_39_54, n_39_53, n_39_52, n_39_51, n_39_50, 
    n_39_49, n_39_48, n_39_47, n_39_46, n_39_45, n_39_44, n_39_43, n_39_42, n_39_41, 
    n_39_40, n_39_39, n_39_38, n_39_37, n_39_36, n_39_35, n_39_34, n_39_33, n_39_32, 
    uc_6}), .b ({\c1[2][31] , \c1[2][30] , \c1[2][29] , \c1[2][28] , \c1[2][27] , 
    \c1[2][26] , \c1[2][25] , \c1[2][24] , \c1[2][23] , \c1[2][22] , \c1[2][21] , 
    \c1[2][20] , \c1[2][19] , \c1[2][18] , \c1[2][17] , \c1[2][16] , \c1[2][15] , 
    \c1[2][14] , \c1[2][13] , \c1[2][12] , \c1[2][11] , \c1[2][10] , \c1[2][9] , 
    \c1[2][8] , \c1[2][7] , \c1[2][6] , \c1[2][5] , \c1[2][4] , \c1[2][3] , \c1[2][2] , 
    \c1[2][1] , \c1[2][0] }), .c ({uc_7, \partial_reg[5][30] , \partial_reg[5][29] , 
    \partial_reg[5][28] , \partial_reg[5][27] , \partial_reg[5][26] , \partial_reg[5][25] , 
    \partial_reg[5][24] , \partial_reg[5][23] , \partial_reg[5][22] , \partial_reg[5][21] , 
    \partial_reg[5][20] , \partial_reg[5][19] , \partial_reg[5][18] , \partial_reg[5][17] , 
    \partial_reg[5][16] , \partial_reg[5][15] , \partial_reg[5][14] , \partial_reg[5][13] , 
    \partial_reg[5][12] , \partial_reg[5][11] , \partial_reg[5][10] , \partial_reg[5][9] , 
    \partial_reg[5][8] , \partial_reg[5][7] , \partial_reg[5][6] , \partial_reg[5][5] , 
    \partial_reg[5][4] , \partial_reg[5][3] , \partial_reg[5][2] , \partial_reg[5][1] , 
    \partial_reg[5][0] }));
PartialAdder__1_283 genblk1_2_p2 (.c1 ({\c1[2][31] , \c1[2][30] , \c1[2][29] , \c1[2][28] , 
    \c1[2][27] , \c1[2][26] , \c1[2][25] , \c1[2][24] , \c1[2][23] , \c1[2][22] , 
    \c1[2][21] , \c1[2][20] , \c1[2][19] , \c1[2][18] , \c1[2][17] , \c1[2][16] , 
    \c1[2][15] , \c1[2][14] , \c1[2][13] , \c1[2][12] , \c1[2][11] , \c1[2][10] , 
    \c1[2][9] , \c1[2][8] , \c1[2][7] , \c1[2][6] , \c1[2][5] , \c1[2][4] , \c1[2][3] , 
    \c1[2][2] , \c1[2][1] , \c1[2][0] }), .s1 ({uc_5, n_39_62, n_39_61, n_39_60, 
    n_39_59, n_39_58, n_39_57, n_39_56, n_39_55, n_39_54, n_39_53, n_39_52, n_39_51, 
    n_39_50, n_39_49, n_39_48, n_39_47, n_39_46, n_39_45, n_39_44, n_39_43, n_39_42, 
    n_39_41, n_39_40, n_39_39, n_39_38, n_39_37, n_39_36, n_39_35, n_39_34, n_39_33, 
    n_39_32, n_1}), .a ({\partial_reg[3][31] , n_39_30, n_39_29, n_39_28, n_39_27, 
    n_39_26, n_39_25, n_39_24, n_39_23, n_39_22, n_39_21, n_39_20, n_39_19, n_39_18, 
    n_39_17, n_39_16, n_39_15, n_39_14, n_39_13, n_39_12, n_39_11, n_39_10, n_39_9, 
    n_39_8, n_39_7, n_39_6, n_39_5, n_39_4, n_39_3, n_39_2, n_39_1, n_39_0, uc_3})
    , .b ({\c1[1][31] , \c1[1][30] , \c1[1][29] , \c1[1][28] , \c1[1][27] , \c1[1][26] , 
    \c1[1][25] , \c1[1][24] , \c1[1][23] , \c1[1][22] , \c1[1][21] , \c1[1][20] , 
    \c1[1][19] , \c1[1][18] , \c1[1][17] , \c1[1][16] , \c1[1][15] , \c1[1][14] , 
    \c1[1][13] , \c1[1][12] , \c1[1][11] , \c1[1][10] , \c1[1][9] , \c1[1][8] , \c1[1][7] , 
    \c1[1][6] , \c1[1][5] , \c1[1][4] , \c1[1][3] , \c1[1][2] , \c1[1][1] , \c1[1][0] })
    , .c ({uc_4, \partial_reg[4][30] , \partial_reg[4][29] , \partial_reg[4][28] , 
    \partial_reg[4][27] , \partial_reg[4][26] , \partial_reg[4][25] , \partial_reg[4][24] , 
    \partial_reg[4][23] , \partial_reg[4][22] , \partial_reg[4][21] , \partial_reg[4][20] , 
    \partial_reg[4][19] , \partial_reg[4][18] , \partial_reg[4][17] , \partial_reg[4][16] , 
    \partial_reg[4][15] , \partial_reg[4][14] , \partial_reg[4][13] , \partial_reg[4][12] , 
    \partial_reg[4][11] , \partial_reg[4][10] , \partial_reg[4][9] , \partial_reg[4][8] , 
    \partial_reg[4][7] , \partial_reg[4][6] , \partial_reg[4][5] , \partial_reg[4][4] , 
    \partial_reg[4][3] , \partial_reg[4][2] , \partial_reg[4][1] , \partial_reg[4][0] }));
PartialAdder__1_186 genblk1_1_p2 (.c1 ({\c1[1][31] , \c1[1][30] , \c1[1][29] , \c1[1][28] , 
    \c1[1][27] , \c1[1][26] , \c1[1][25] , \c1[1][24] , \c1[1][23] , \c1[1][22] , 
    \c1[1][21] , \c1[1][20] , \c1[1][19] , \c1[1][18] , \c1[1][17] , \c1[1][16] , 
    \c1[1][15] , \c1[1][14] , \c1[1][13] , \c1[1][12] , \c1[1][11] , \c1[1][10] , 
    \c1[1][9] , \c1[1][8] , \c1[1][7] , \c1[1][6] , \c1[1][5] , \c1[1][4] , \c1[1][3] , 
    \c1[1][2] , \c1[1][1] , \c1[1][0] }), .s1 ({uc_2, n_39_30, n_39_29, n_39_28, 
    n_39_27, n_39_26, n_39_25, n_39_24, n_39_23, n_39_22, n_39_21, n_39_20, n_39_19, 
    n_39_18, n_39_17, n_39_16, n_39_15, n_39_14, n_39_13, n_39_12, n_39_11, n_39_10, 
    n_39_9, n_39_8, n_39_7, n_39_6, n_39_5, n_39_4, n_39_3, n_39_2, n_39_1, n_39_0, 
    n_0}), .a ({\partial_reg[2][31] , \s1[0][31] , \s1[0][30] , \s1[0][29] , \s1[0][28] , 
    \s1[0][27] , \s1[0][26] , \s1[0][25] , \s1[0][24] , \s1[0][23] , \s1[0][22] , 
    \s1[0][21] , \s1[0][20] , \s1[0][19] , \s1[0][18] , \s1[0][17] , \s1[0][16] , 
    \s1[0][15] , \s1[0][14] , \s1[0][13] , \s1[0][12] , \s1[0][11] , \s1[0][10] , 
    \s1[0][9] , \s1[0][8] , \s1[0][7] , \s1[0][6] , \s1[0][5] , \s1[0][4] , \s1[0][3] , 
    \s1[0][2] , \s1[0][1] , uc_0}), .b ({\c1[0][31] , \c1[0][30] , \c1[0][29] , \c1[0][28] , 
    \c1[0][27] , \c1[0][26] , \c1[0][25] , \c1[0][24] , \c1[0][23] , \c1[0][22] , 
    \c1[0][21] , \c1[0][20] , \c1[0][19] , \c1[0][18] , \c1[0][17] , \c1[0][16] , 
    \c1[0][15] , \c1[0][14] , \c1[0][13] , \c1[0][12] , \c1[0][11] , \c1[0][10] , 
    \c1[0][9] , \c1[0][8] , \c1[0][7] , \c1[0][6] , \c1[0][5] , \c1[0][4] , \c1[0][3] , 
    \c1[0][2] , \c1[0][1] , \c1[0][0] }), .c ({uc_1, \partial_reg[3][30] , \partial_reg[3][29] , 
    \partial_reg[3][28] , \partial_reg[3][27] , \partial_reg[3][26] , \partial_reg[3][25] , 
    \partial_reg[3][24] , \partial_reg[3][23] , \partial_reg[3][22] , \partial_reg[3][21] , 
    \partial_reg[3][20] , \partial_reg[3][19] , \partial_reg[3][18] , \partial_reg[3][17] , 
    \partial_reg[3][16] , \partial_reg[3][15] , \partial_reg[3][14] , \partial_reg[3][13] , 
    \partial_reg[3][12] , \partial_reg[3][11] , \partial_reg[3][10] , \partial_reg[3][9] , 
    \partial_reg[3][8] , \partial_reg[3][7] , \partial_reg[3][6] , \partial_reg[3][5] , 
    \partial_reg[3][4] , \partial_reg[3][3] , \partial_reg[3][2] , \partial_reg[3][1] , 
    \partial_reg[3][0] }));

endmodule //TreeMultiplierCirc

module TreeMultiplier (a, b, clk, data);

output [63:0] data;
input [31:0] a;
input [31:0] b;
input clk;
wire \out[63] ;
wire \out[62] ;
wire \out[61] ;
wire \out[60] ;
wire \out[59] ;
wire \out[58] ;
wire \out[57] ;
wire \out[56] ;
wire \out[55] ;
wire \out[54] ;
wire \out[53] ;
wire \out[52] ;
wire \out[51] ;
wire \out[50] ;
wire \out[49] ;
wire \out[48] ;
wire \out[47] ;
wire \out[46] ;
wire \out[45] ;
wire \out[44] ;
wire \out[43] ;
wire \out[42] ;
wire \out[41] ;
wire \out[40] ;
wire \out[39] ;
wire \out[38] ;
wire \out[37] ;
wire \out[36] ;
wire \out[35] ;
wire \out[34] ;
wire \out[33] ;
wire \out[32] ;
wire \out[31] ;
wire \out[30] ;
wire \out[29] ;
wire \out[28] ;
wire \out[27] ;
wire \out[26] ;
wire \out[25] ;
wire \out[24] ;
wire \out[23] ;
wire \out[22] ;
wire \out[21] ;
wire \out[20] ;
wire \out[19] ;
wire \out[18] ;
wire \out[17] ;
wire \out[16] ;
wire \out[15] ;
wire \out[14] ;
wire \out[13] ;
wire \out[12] ;
wire \out[11] ;
wire \out[10] ;
wire \out[9] ;
wire \out[8] ;
wire \out[7] ;
wire \out[6] ;
wire \out[5] ;
wire \out[4] ;
wire \out[3] ;
wire \out[2] ;
wire \out[1] ;
wire \out[0] ;
wire \c[31] ;
wire \c[30] ;
wire \c[29] ;
wire \c[28] ;
wire \c[27] ;
wire \c[26] ;
wire \c[25] ;
wire \c[24] ;
wire \c[23] ;
wire \c[22] ;
wire \c[21] ;
wire \c[20] ;
wire \c[19] ;
wire \c[18] ;
wire \c[17] ;
wire \c[16] ;
wire \c[15] ;
wire \c[14] ;
wire \c[13] ;
wire \c[12] ;
wire \c[11] ;
wire \c[10] ;
wire \c[9] ;
wire \c[8] ;
wire \c[7] ;
wire \c[6] ;
wire \c[5] ;
wire \c[4] ;
wire \c[3] ;
wire \c[2] ;
wire \c[1] ;
wire \c[0] ;
wire \d[31] ;
wire \d[30] ;
wire \d[29] ;
wire \d[28] ;
wire \d[27] ;
wire \d[26] ;
wire \d[25] ;
wire \d[24] ;
wire \d[23] ;
wire \d[22] ;
wire \d[21] ;
wire \d[20] ;
wire \d[19] ;
wire \d[18] ;
wire \d[17] ;
wire \d[16] ;
wire \d[15] ;
wire \d[14] ;
wire \d[13] ;
wire \d[12] ;
wire \d[11] ;
wire \d[10] ;
wire \d[9] ;
wire \d[8] ;
wire \d[7] ;
wire \d[6] ;
wire \d[5] ;
wire \d[4] ;
wire \d[3] ;
wire \d[2] ;
wire \d[1] ;
wire \d[0] ;
wire CTS_n83;
wire CTS_n181;
wire CTS_n207;
wire CLOCK_n340;


Register__parameterized0 Register_inst3 (.out ({data[63], data[62], data[61], data[60], 
    data[59], data[58], data[57], data[56], data[55], data[54], data[53], data[52], 
    data[51], data[50], data[49], data[48], data[47], data[46], data[45], data[44], 
    data[43], data[42], data[41], data[40], data[39], data[38], data[37], data[36], 
    data[35], data[34], data[33], data[32], data[31], data[30], data[29], data[28], 
    data[27], data[26], data[25], data[24], data[23], data[22], data[21], data[20], 
    data[19], data[18], data[17], data[16], data[15], data[14], data[13], data[12], 
    data[11], data[10], data[9], data[8], data[7], data[6], data[5], data[4], data[3], 
    data[2], data[1], data[0]}), .in ({\out[63] , \out[62] , \out[61] , \out[60] , 
    \out[59] , \out[58] , \out[57] , \out[56] , \out[55] , \out[54] , \out[53] , 
    \out[52] , \out[51] , \out[50] , \out[49] , \out[48] , \out[47] , \out[46] , 
    \out[45] , \out[44] , \out[43] , \out[42] , \out[41] , \out[40] , \out[39] , 
    \out[38] , \out[37] , \out[36] , \out[35] , \out[34] , \out[33] , \out[32] , 
    \out[31] , \out[30] , \out[29] , \out[28] , \out[27] , \out[26] , \out[25] , 
    \out[24] , \out[23] , \out[22] , \out[21] , \out[20] , \out[19] , \out[18] , 
    \out[17] , \out[16] , \out[15] , \out[14] , \out[13] , \out[12] , \out[11] , 
    \out[10] , \out[9] , \out[8] , \out[7] , \out[6] , \out[5] , \out[4] , \out[3] , 
    \out[2] , \out[1] , \out[0] }), .clk_CTSPP_21 (CTS_n83), .clk_CTSPP_62 (CTS_n207)
    , .clk_CTSPP_72 (CLOCK_n340));
Register Register_inst2 (.out ({\d[31] , \d[30] , \d[29] , \d[28] , \d[27] , \d[26] , 
    \d[25] , \d[24] , \d[23] , \d[22] , \d[21] , \d[20] , \d[19] , \d[18] , \d[17] , 
    \d[16] , \d[15] , \d[14] , \d[13] , \d[12] , \d[11] , \d[10] , \d[9] , \d[8] , 
    \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , \d[2] , \d[1] , \d[0] }), .clk_CTSPP_48 (CTS_n181)
    , .clk_CTSPP_61 (CTS_n207), .in ({b[31], b[30], b[29], b[28], b[27], b[26], b[25], 
    b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], b[15], b[14], 
    b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], 
    b[0]}), .clk_CTSPP_70 (CLOCK_n340));
Register__5_0 Register_inst1 (.out ({\c[31] , \c[30] , \c[29] , \c[28] , \c[27] , 
    \c[26] , \c[25] , \c[24] , \c[23] , \c[22] , \c[21] , \c[20] , \c[19] , \c[18] , 
    \c[17] , \c[16] , \c[15] , \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , 
    \c[8] , \c[7] , \c[6] , \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] }), .clk_CTSPP_23 (CTS_n83)
    , .in ({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], 
    a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], 
    a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), .clk_CTSPP_52 (CTS_n181)
    , .clk_CTSPP_60 (CLOCK_n340));
TreeMultiplierCirc t1 (.out ({\out[63] , \out[62] , \out[61] , \out[60] , \out[59] , 
    \out[58] , \out[57] , \out[56] , \out[55] , \out[54] , \out[53] , \out[52] , 
    \out[51] , \out[50] , \out[49] , \out[48] , \out[47] , \out[46] , \out[45] , 
    \out[44] , \out[43] , \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , 
    \out[37] , \out[36] , \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , 
    \out[30] , \out[29] , \out[28] , \out[27] , \out[26] , \out[25] , \out[24] , 
    \out[23] , \out[22] , \out[21] , \out[20] , \out[19] , \out[18] , \out[17] , 
    \out[16] , \out[15] , \out[14] , \out[13] , \out[12] , \out[11] , \out[10] , 
    \out[9] , \out[8] , \out[7] , \out[6] , \out[5] , \out[4] , \out[3] , \out[2] , 
    \out[1] , \out[0] }), .a ({\c[31] , \c[30] , \c[29] , \c[28] , \c[27] , \c[26] , 
    \c[25] , \c[24] , \c[23] , \c[22] , \c[21] , \c[20] , \c[19] , \c[18] , \c[17] , 
    \c[16] , \c[15] , \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , \c[8] , 
    \c[7] , \c[6] , \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] }), .b ({\d[31] , 
    \d[30] , \d[29] , \d[28] , \d[27] , \d[26] , \d[25] , \d[24] , \d[23] , \d[22] , 
    \d[21] , \d[20] , \d[19] , \d[18] , \d[17] , \d[16] , \d[15] , \d[14] , \d[13] , 
    \d[12] , \d[11] , \d[10] , \d[9] , \d[8] , \d[7] , \d[6] , \d[5] , \d[4] , \d[3] , 
    \d[2] , \d[1] , \d[0] }));
CLKBUF_X2 CTS_L1_c1_c45 (.Z (CLOCK_n340), .A (clk));

endmodule //TreeMultiplier


