/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Oct 31 17:17:33 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 686356441 */

module halfAdder__0_12(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_13(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_12 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_17(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
endmodule

module fullAdder__0_21(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_17 h2 (.x(y), .y(cin), .sum(sum), .cout());
endmodule

module halfAdder__0_28(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_29(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_28 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_36(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_37(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_36 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_44(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_45(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_44 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_52(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_53(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_52 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_60(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_61(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_60 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_68(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_69(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_68 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_76(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_77(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_76 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_84(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_85(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_84 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_92(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_93(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_92 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_100(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_101(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_100 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_108(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_109(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_108 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_116(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_117(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_116 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_124(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_125(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_124 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_132(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_133(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_132 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_140(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_141(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_140 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_148(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_149(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_148 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_156(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_157(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_156 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_164(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_165(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_164 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_172(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_173(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_172 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_180(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_181(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_180 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_188(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_189(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_188 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_196(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_197(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_196 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_204(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_205(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_204 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_212(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_212 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_220(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_221(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_220 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_228(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_229(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_228 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_236(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_237(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_236 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_244(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_245(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_244 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_252(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_253(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_252 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_260(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_261(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_260 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_268(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_269(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_268 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_276(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_277(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   halfAdder__0_276 h1 (.x(x), .y(y), .sum(sum), .cout(cout));
endmodule

module halfAdder__0_284(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_281(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_285(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_284 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_281 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_292(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_289(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_293(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_292 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_289 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_300(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_297(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_301(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_300 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_297 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_308(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_305(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_309(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_308 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_305 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_316(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_313(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_317(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_316 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_313 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_324(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_321(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_325(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_324 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_321 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_332(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_329(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_333(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_332 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_329 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_340(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_337(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_341(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_340 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_337 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_348(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_345(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_349(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_348 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_345 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_356(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_353(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_357(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_356 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_353 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_364(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_361(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_365(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_364 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_361 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_372(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_369(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_373(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_372 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_369 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_380(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_377(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_381(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_380 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_377 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_388(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_385(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_389(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_388 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_385 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_396(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_393(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_397(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_396 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_393 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_404(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_401(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_405(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_404 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_401 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_412(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_409(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_413(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_412 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_409 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_420(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_417(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_421(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_420 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_417 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_428(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_425(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_429(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_428 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_425 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_436(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_433(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_437(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_436 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_433 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_444(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_441(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_445(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_444 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_441 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_452(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_449(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_453(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_452 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_449 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_460(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_457(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_461(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_460 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_457 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_468(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_465(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_469(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_468 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_465 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_476(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_473(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_477(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_476 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_473 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_484(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_481(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_485(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_484 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_481 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_492(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_489(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_493(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_492 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_489 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_500(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_497(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_501(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_500 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_497 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_508(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder__0_505(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder__0_509(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_508 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder__0_505 h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module halfAdder__0_5(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module halfAdder(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module fullAdder(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire halfCarry1;
   wire halfSum;
   wire halfCarry2;

   halfAdder__0_5 h1 (.x(x), .y(y), .sum(halfSum), .cout(halfCarry1));
   halfAdder h2 (.x(halfSum), .y(cin), .sum(sum), .cout(halfCarry2));
   OR2_X1 i_0_0 (.A1(halfCarry2), .A2(halfCarry1), .ZN(cout));
endmodule

module carrySaveAdder(a, b, cin, sum, cout);
   input [31:0]a;
   input [31:0]b;
   input cin;
   output [31:0]sum;
   output cout;

   wire [30:0]halfcarry;
   wire [31:0]halfcout;
   wire [31:0]halfsum;

   fullAdder__0_13 fulladder_f2 (.x(halfsum[1]), .y(halfcout[0]), .cin(), 
      .sum(sum[1]), .cout(halfcarry[0]));
   fullAdder__0_21 fulladder_f3 (.x(), .y(halfcout[31]), .cin(halfcarry[30]), 
      .sum(cout), .cout());
   fullAdder__0_29 genblk1_0_fulladder_f1 (.x(a[0]), .y(b[0]), .cin(), .sum(
      sum[0]), .cout(halfcout[0]));
   fullAdder__0_37 genblk1_1_fulladder_f1 (.x(a[1]), .y(b[1]), .cin(), .sum(
      halfsum[1]), .cout(halfcout[1]));
   fullAdder__0_45 genblk1_2_fulladder_f1 (.x(a[2]), .y(b[2]), .cin(), .sum(
      halfsum[2]), .cout(halfcout[2]));
   fullAdder__0_53 genblk1_3_fulladder_f1 (.x(a[3]), .y(b[3]), .cin(), .sum(
      halfsum[3]), .cout(halfcout[3]));
   fullAdder__0_61 genblk1_4_fulladder_f1 (.x(a[4]), .y(b[4]), .cin(), .sum(
      halfsum[4]), .cout(halfcout[4]));
   fullAdder__0_69 genblk1_5_fulladder_f1 (.x(a[5]), .y(b[5]), .cin(), .sum(
      halfsum[5]), .cout(halfcout[5]));
   fullAdder__0_77 genblk1_6_fulladder_f1 (.x(a[6]), .y(b[6]), .cin(), .sum(
      halfsum[6]), .cout(halfcout[6]));
   fullAdder__0_85 genblk1_7_fulladder_f1 (.x(a[7]), .y(b[7]), .cin(), .sum(
      halfsum[7]), .cout(halfcout[7]));
   fullAdder__0_93 genblk1_8_fulladder_f1 (.x(a[8]), .y(b[8]), .cin(), .sum(
      halfsum[8]), .cout(halfcout[8]));
   fullAdder__0_101 genblk1_9_fulladder_f1 (.x(a[9]), .y(b[9]), .cin(), .sum(
      halfsum[9]), .cout(halfcout[9]));
   fullAdder__0_109 genblk1_10_fulladder_f1 (.x(a[10]), .y(b[10]), .cin(), 
      .sum(halfsum[10]), .cout(halfcout[10]));
   fullAdder__0_117 genblk1_11_fulladder_f1 (.x(a[11]), .y(b[11]), .cin(), 
      .sum(halfsum[11]), .cout(halfcout[11]));
   fullAdder__0_125 genblk1_12_fulladder_f1 (.x(a[12]), .y(b[12]), .cin(), 
      .sum(halfsum[12]), .cout(halfcout[12]));
   fullAdder__0_133 genblk1_13_fulladder_f1 (.x(a[13]), .y(b[13]), .cin(), 
      .sum(halfsum[13]), .cout(halfcout[13]));
   fullAdder__0_141 genblk1_14_fulladder_f1 (.x(a[14]), .y(b[14]), .cin(), 
      .sum(halfsum[14]), .cout(halfcout[14]));
   fullAdder__0_149 genblk1_15_fulladder_f1 (.x(a[15]), .y(b[15]), .cin(), 
      .sum(halfsum[15]), .cout(halfcout[15]));
   fullAdder__0_157 genblk1_16_fulladder_f1 (.x(a[16]), .y(b[16]), .cin(), 
      .sum(halfsum[16]), .cout(halfcout[16]));
   fullAdder__0_165 genblk1_17_fulladder_f1 (.x(a[17]), .y(b[17]), .cin(), 
      .sum(halfsum[17]), .cout(halfcout[17]));
   fullAdder__0_173 genblk1_18_fulladder_f1 (.x(a[18]), .y(b[18]), .cin(), 
      .sum(halfsum[18]), .cout(halfcout[18]));
   fullAdder__0_181 genblk1_19_fulladder_f1 (.x(a[19]), .y(b[19]), .cin(), 
      .sum(halfsum[19]), .cout(halfcout[19]));
   fullAdder__0_189 genblk1_20_fulladder_f1 (.x(a[20]), .y(b[20]), .cin(), 
      .sum(halfsum[20]), .cout(halfcout[20]));
   fullAdder__0_197 genblk1_21_fulladder_f1 (.x(a[21]), .y(b[21]), .cin(), 
      .sum(halfsum[21]), .cout(halfcout[21]));
   fullAdder__0_205 genblk1_22_fulladder_f1 (.x(a[22]), .y(b[22]), .cin(), 
      .sum(halfsum[22]), .cout(halfcout[22]));
   fullAdder__0_213 genblk1_23_fulladder_f1 (.x(a[23]), .y(b[23]), .cin(), 
      .sum(halfsum[23]), .cout(halfcout[23]));
   fullAdder__0_221 genblk1_24_fulladder_f1 (.x(a[24]), .y(b[24]), .cin(), 
      .sum(halfsum[24]), .cout(halfcout[24]));
   fullAdder__0_229 genblk1_25_fulladder_f1 (.x(a[25]), .y(b[25]), .cin(), 
      .sum(halfsum[25]), .cout(halfcout[25]));
   fullAdder__0_237 genblk1_26_fulladder_f1 (.x(a[26]), .y(b[26]), .cin(), 
      .sum(halfsum[26]), .cout(halfcout[26]));
   fullAdder__0_245 genblk1_27_fulladder_f1 (.x(a[27]), .y(b[27]), .cin(), 
      .sum(halfsum[27]), .cout(halfcout[27]));
   fullAdder__0_253 genblk1_28_fulladder_f1 (.x(a[28]), .y(b[28]), .cin(), 
      .sum(halfsum[28]), .cout(halfcout[28]));
   fullAdder__0_261 genblk1_29_fulladder_f1 (.x(a[29]), .y(b[29]), .cin(), 
      .sum(halfsum[29]), .cout(halfcout[29]));
   fullAdder__0_269 genblk1_30_fulladder_f1 (.x(a[30]), .y(b[30]), .cin(), 
      .sum(halfsum[30]), .cout(halfcout[30]));
   fullAdder__0_277 genblk1_31_fulladder_f1 (.x(a[31]), .y(b[31]), .cin(), 
      .sum(halfsum[31]), .cout(halfcout[31]));
   fullAdder__0_285 genblk2_1_f3 (.x(halfsum[2]), .y(halfcout[1]), .cin(
      halfcarry[0]), .sum(sum[2]), .cout(halfcarry[1]));
   fullAdder__0_293 genblk2_2_f3 (.x(halfsum[3]), .y(halfcout[2]), .cin(
      halfcarry[1]), .sum(sum[3]), .cout(halfcarry[2]));
   fullAdder__0_301 genblk2_3_f3 (.x(halfsum[4]), .y(halfcout[3]), .cin(
      halfcarry[2]), .sum(sum[4]), .cout(halfcarry[3]));
   fullAdder__0_309 genblk2_4_f3 (.x(halfsum[5]), .y(halfcout[4]), .cin(
      halfcarry[3]), .sum(sum[5]), .cout(halfcarry[4]));
   fullAdder__0_317 genblk2_5_f3 (.x(halfsum[6]), .y(halfcout[5]), .cin(
      halfcarry[4]), .sum(sum[6]), .cout(halfcarry[5]));
   fullAdder__0_325 genblk2_6_f3 (.x(halfsum[7]), .y(halfcout[6]), .cin(
      halfcarry[5]), .sum(sum[7]), .cout(halfcarry[6]));
   fullAdder__0_333 genblk2_7_f3 (.x(halfsum[8]), .y(halfcout[7]), .cin(
      halfcarry[6]), .sum(sum[8]), .cout(halfcarry[7]));
   fullAdder__0_341 genblk2_8_f3 (.x(halfsum[9]), .y(halfcout[8]), .cin(
      halfcarry[7]), .sum(sum[9]), .cout(halfcarry[8]));
   fullAdder__0_349 genblk2_9_f3 (.x(halfsum[10]), .y(halfcout[9]), .cin(
      halfcarry[8]), .sum(sum[10]), .cout(halfcarry[9]));
   fullAdder__0_357 genblk2_10_f3 (.x(halfsum[11]), .y(halfcout[10]), .cin(
      halfcarry[9]), .sum(sum[11]), .cout(halfcarry[10]));
   fullAdder__0_365 genblk2_11_f3 (.x(halfsum[12]), .y(halfcout[11]), .cin(
      halfcarry[10]), .sum(sum[12]), .cout(halfcarry[11]));
   fullAdder__0_373 genblk2_12_f3 (.x(halfsum[13]), .y(halfcout[12]), .cin(
      halfcarry[11]), .sum(sum[13]), .cout(halfcarry[12]));
   fullAdder__0_381 genblk2_13_f3 (.x(halfsum[14]), .y(halfcout[13]), .cin(
      halfcarry[12]), .sum(sum[14]), .cout(halfcarry[13]));
   fullAdder__0_389 genblk2_14_f3 (.x(halfsum[15]), .y(halfcout[14]), .cin(
      halfcarry[13]), .sum(sum[15]), .cout(halfcarry[14]));
   fullAdder__0_397 genblk2_15_f3 (.x(halfsum[16]), .y(halfcout[15]), .cin(
      halfcarry[14]), .sum(sum[16]), .cout(halfcarry[15]));
   fullAdder__0_405 genblk2_16_f3 (.x(halfsum[17]), .y(halfcout[16]), .cin(
      halfcarry[15]), .sum(sum[17]), .cout(halfcarry[16]));
   fullAdder__0_413 genblk2_17_f3 (.x(halfsum[18]), .y(halfcout[17]), .cin(
      halfcarry[16]), .sum(sum[18]), .cout(halfcarry[17]));
   fullAdder__0_421 genblk2_18_f3 (.x(halfsum[19]), .y(halfcout[18]), .cin(
      halfcarry[17]), .sum(sum[19]), .cout(halfcarry[18]));
   fullAdder__0_429 genblk2_19_f3 (.x(halfsum[20]), .y(halfcout[19]), .cin(
      halfcarry[18]), .sum(sum[20]), .cout(halfcarry[19]));
   fullAdder__0_437 genblk2_20_f3 (.x(halfsum[21]), .y(halfcout[20]), .cin(
      halfcarry[19]), .sum(sum[21]), .cout(halfcarry[20]));
   fullAdder__0_445 genblk2_21_f3 (.x(halfsum[22]), .y(halfcout[21]), .cin(
      halfcarry[20]), .sum(sum[22]), .cout(halfcarry[21]));
   fullAdder__0_453 genblk2_22_f3 (.x(halfsum[23]), .y(halfcout[22]), .cin(
      halfcarry[21]), .sum(sum[23]), .cout(halfcarry[22]));
   fullAdder__0_461 genblk2_23_f3 (.x(halfsum[24]), .y(halfcout[23]), .cin(
      halfcarry[22]), .sum(sum[24]), .cout(halfcarry[23]));
   fullAdder__0_469 genblk2_24_f3 (.x(halfsum[25]), .y(halfcout[24]), .cin(
      halfcarry[23]), .sum(sum[25]), .cout(halfcarry[24]));
   fullAdder__0_477 genblk2_25_f3 (.x(halfsum[26]), .y(halfcout[25]), .cin(
      halfcarry[24]), .sum(sum[26]), .cout(halfcarry[25]));
   fullAdder__0_485 genblk2_26_f3 (.x(halfsum[27]), .y(halfcout[26]), .cin(
      halfcarry[25]), .sum(sum[27]), .cout(halfcarry[26]));
   fullAdder__0_493 genblk2_27_f3 (.x(halfsum[28]), .y(halfcout[27]), .cin(
      halfcarry[26]), .sum(sum[28]), .cout(halfcarry[27]));
   fullAdder__0_501 genblk2_28_f3 (.x(halfsum[29]), .y(halfcout[28]), .cin(
      halfcarry[27]), .sum(sum[29]), .cout(halfcarry[28]));
   fullAdder__0_509 genblk2_29_f3 (.x(halfsum[30]), .y(halfcout[29]), .cin(
      halfcarry[28]), .sum(sum[30]), .cout(halfcarry[29]));
   fullAdder genblk2_30_f3 (.x(halfsum[31]), .y(halfcout[30]), .cin(
      halfcarry[29]), .sum(sum[31]), .cout(halfcarry[30]));
endmodule
