
// 	Wed Jan  4 04:39:12 2023
//	vlsi
//	localhost.localdomain

module datapath__0_29 (input_plus, inputM_inv22, inputM);

output [31:0] inputM_inv22;
input [31:0] inputM;
input input_plus;
wire n_40;
wire n_0;
wire n_43;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_32;
wire n_30;
wire n_29;
wire n_27;
wire n_26;
wire n_24;
wire n_23;
wire n_21;
wire n_20;
wire n_18;
wire n_17;
wire n_15;
wire n_14;
wire n_12;
wire n_11;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_1;
wire n_2;
wire n_5;
wire n_4;
wire n_3;
wire n_42;
wire n_41;
wire n_10;
wire n_13;
wire n_16;
wire n_19;
wire n_22;
wire n_25;
wire n_28;
wire n_31;
wire n_33;


INV_X1 i_75 (.ZN (n_43), .A (input_plus));
INV_X1 i_74 (.ZN (n_42), .A (inputM[28]));
INV_X1 i_73 (.ZN (n_41), .A (inputM[25]));
OR3_X1 i_72 (.ZN (n_40), .A1 (n_43), .A2 (inputM[1]), .A3 (inputM[0]));
OR2_X1 i_71 (.ZN (n_39), .A1 (n_40), .A2 (inputM[2]));
OR2_X1 i_70 (.ZN (n_38), .A1 (n_39), .A2 (inputM[3]));
OR2_X1 i_69 (.ZN (n_37), .A1 (n_38), .A2 (inputM[4]));
NOR2_X1 i_68 (.ZN (n_36), .A1 (n_37), .A2 (inputM[5]));
NOR3_X1 i_67 (.ZN (n_35), .A1 (n_37), .A2 (inputM[5]), .A3 (inputM[6]));
NOR4_X1 i_66 (.ZN (n_34), .A1 (n_37), .A2 (inputM[5]), .A3 (inputM[6]), .A4 (inputM[7]));
INV_X1 i_65 (.ZN (n_33), .A (n_34));
NOR2_X1 i_64 (.ZN (n_32), .A1 (n_33), .A2 (inputM[8]));
INV_X1 i_63 (.ZN (n_31), .A (n_32));
NOR2_X1 i_62 (.ZN (n_30), .A1 (n_31), .A2 (inputM[9]));
NOR3_X1 i_61 (.ZN (n_29), .A1 (n_31), .A2 (inputM[9]), .A3 (inputM[10]));
INV_X1 i_60 (.ZN (n_28), .A (n_29));
NOR2_X1 i_59 (.ZN (n_27), .A1 (n_28), .A2 (inputM[11]));
NOR3_X1 i_58 (.ZN (n_26), .A1 (n_28), .A2 (inputM[11]), .A3 (inputM[12]));
INV_X1 i_57 (.ZN (n_25), .A (n_26));
NOR2_X1 i_56 (.ZN (n_24), .A1 (n_25), .A2 (inputM[13]));
NOR3_X1 i_55 (.ZN (n_23), .A1 (n_25), .A2 (inputM[13]), .A3 (inputM[14]));
INV_X1 i_54 (.ZN (n_22), .A (n_23));
NOR2_X1 i_53 (.ZN (n_21), .A1 (n_22), .A2 (inputM[15]));
NOR3_X1 i_52 (.ZN (n_20), .A1 (n_22), .A2 (inputM[15]), .A3 (inputM[16]));
INV_X1 i_51 (.ZN (n_19), .A (n_20));
NOR2_X1 i_50 (.ZN (n_18), .A1 (n_19), .A2 (inputM[17]));
NOR3_X1 i_49 (.ZN (n_17), .A1 (n_19), .A2 (inputM[17]), .A3 (inputM[18]));
INV_X1 i_48 (.ZN (n_16), .A (n_17));
NOR2_X1 i_47 (.ZN (n_15), .A1 (n_16), .A2 (inputM[19]));
NOR3_X1 i_46 (.ZN (n_14), .A1 (n_16), .A2 (inputM[19]), .A3 (inputM[20]));
INV_X1 i_45 (.ZN (n_13), .A (n_14));
NOR2_X1 i_44 (.ZN (n_12), .A1 (n_13), .A2 (inputM[21]));
NOR3_X1 i_43 (.ZN (n_11), .A1 (n_13), .A2 (inputM[21]), .A3 (inputM[22]));
INV_X1 i_42 (.ZN (n_10), .A (n_11));
NOR2_X1 i_41 (.ZN (n_9), .A1 (n_10), .A2 (inputM[23]));
NOR3_X1 i_40 (.ZN (n_8), .A1 (n_10), .A2 (inputM[23]), .A3 (inputM[24]));
NAND2_X1 i_39 (.ZN (n_7), .A1 (n_8), .A2 (n_41));
NOR3_X1 i_38 (.ZN (n_6), .A1 (n_7), .A2 (inputM[26]), .A3 (inputM[27]));
NAND2_X1 i_37 (.ZN (n_5), .A1 (n_6), .A2 (n_42));
NOR2_X1 i_36 (.ZN (n_4), .A1 (n_5), .A2 (inputM[29]));
NOR3_X1 i_35 (.ZN (n_3), .A1 (n_5), .A2 (inputM[29]), .A3 (inputM[30]));
XNOR2_X1 i_34 (.ZN (inputM_inv22[31]), .A (inputM[31]), .B (n_3));
XNOR2_X1 i_33 (.ZN (inputM_inv22[30]), .A (inputM[30]), .B (n_4));
XOR2_X1 i_32 (.Z (inputM_inv22[29]), .A (inputM[29]), .B (n_5));
XNOR2_X1 i_31 (.ZN (inputM_inv22[28]), .A (inputM[28]), .B (n_6));
OAI21_X1 i_30 (.ZN (n_2), .A (inputM[27]), .B1 (n_7), .B2 (inputM[26]));
INV_X1 i_29 (.ZN (n_1), .A (n_2));
NOR2_X1 i_28 (.ZN (inputM_inv22[27]), .A1 (n_6), .A2 (n_1));
XOR2_X1 i_27 (.Z (inputM_inv22[26]), .A (inputM[26]), .B (n_7));
XNOR2_X1 i_26 (.ZN (inputM_inv22[25]), .A (inputM[25]), .B (n_8));
XNOR2_X1 i_25 (.ZN (inputM_inv22[24]), .A (inputM[24]), .B (n_9));
XNOR2_X1 i_24 (.ZN (inputM_inv22[23]), .A (inputM[23]), .B (n_11));
XNOR2_X1 i_23 (.ZN (inputM_inv22[22]), .A (inputM[22]), .B (n_12));
XNOR2_X1 i_22 (.ZN (inputM_inv22[21]), .A (inputM[21]), .B (n_14));
XNOR2_X1 i_21 (.ZN (inputM_inv22[20]), .A (inputM[20]), .B (n_15));
XNOR2_X1 i_20 (.ZN (inputM_inv22[19]), .A (inputM[19]), .B (n_17));
XNOR2_X1 i_19 (.ZN (inputM_inv22[18]), .A (inputM[18]), .B (n_18));
XNOR2_X1 i_18 (.ZN (inputM_inv22[17]), .A (inputM[17]), .B (n_20));
XNOR2_X1 i_17 (.ZN (inputM_inv22[16]), .A (inputM[16]), .B (n_21));
XNOR2_X1 i_16 (.ZN (inputM_inv22[15]), .A (inputM[15]), .B (n_23));
XNOR2_X1 i_15 (.ZN (inputM_inv22[14]), .A (inputM[14]), .B (n_24));
XNOR2_X1 i_14 (.ZN (inputM_inv22[13]), .A (inputM[13]), .B (n_26));
XNOR2_X1 i_13 (.ZN (inputM_inv22[12]), .A (inputM[12]), .B (n_27));
XNOR2_X1 i_12 (.ZN (inputM_inv22[11]), .A (inputM[11]), .B (n_29));
XNOR2_X1 i_11 (.ZN (inputM_inv22[10]), .A (inputM[10]), .B (n_30));
XNOR2_X1 i_10 (.ZN (inputM_inv22[9]), .A (inputM[9]), .B (n_32));
XNOR2_X1 i_9 (.ZN (inputM_inv22[8]), .A (inputM[8]), .B (n_34));
XNOR2_X1 i_8 (.ZN (inputM_inv22[7]), .A (inputM[7]), .B (n_35));
XNOR2_X1 i_7 (.ZN (inputM_inv22[6]), .A (inputM[6]), .B (n_36));
XOR2_X1 i_6 (.Z (inputM_inv22[5]), .A (inputM[5]), .B (n_37));
XOR2_X1 i_5 (.Z (inputM_inv22[4]), .A (inputM[4]), .B (n_38));
XOR2_X1 i_4 (.Z (inputM_inv22[3]), .A (inputM[3]), .B (n_39));
XOR2_X1 i_3 (.Z (inputM_inv22[2]), .A (inputM[2]), .B (n_40));
OAI21_X1 i_2 (.ZN (n_0), .A (inputM[1]), .B1 (n_43), .B2 (inputM[0]));
AND2_X1 i_1 (.ZN (inputM_inv22[1]), .A1 (n_40), .A2 (n_0));
XNOR2_X1 i_0 (.ZN (inputM_inv22[0]), .A (input_plus), .B (inputM[0]));

endmodule //datapath__0_29

module datapath__0_27 (input_plus, inputQ_inv22, inputQ);

output [31:0] inputQ_inv22;
input [31:0] inputQ;
input input_plus;
wire n_40;
wire n_0;
wire n_43;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_32;
wire n_30;
wire n_29;
wire n_27;
wire n_26;
wire n_24;
wire n_23;
wire n_21;
wire n_20;
wire n_18;
wire n_17;
wire n_15;
wire n_14;
wire n_12;
wire n_11;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_1;
wire n_2;
wire n_5;
wire n_4;
wire n_3;
wire n_42;
wire n_41;
wire n_10;
wire n_13;
wire n_16;
wire n_19;
wire n_22;
wire n_25;
wire n_28;
wire n_31;
wire n_33;


INV_X1 i_75 (.ZN (n_43), .A (input_plus));
INV_X1 i_74 (.ZN (n_42), .A (inputQ[28]));
INV_X1 i_73 (.ZN (n_41), .A (inputQ[25]));
OR3_X1 i_72 (.ZN (n_40), .A1 (n_43), .A2 (inputQ[1]), .A3 (inputQ[0]));
OR2_X1 i_71 (.ZN (n_39), .A1 (n_40), .A2 (inputQ[2]));
OR2_X1 i_70 (.ZN (n_38), .A1 (n_39), .A2 (inputQ[3]));
OR2_X1 i_69 (.ZN (n_37), .A1 (n_38), .A2 (inputQ[4]));
NOR2_X1 i_68 (.ZN (n_36), .A1 (n_37), .A2 (inputQ[5]));
NOR3_X1 i_67 (.ZN (n_35), .A1 (n_37), .A2 (inputQ[5]), .A3 (inputQ[6]));
NOR4_X1 i_66 (.ZN (n_34), .A1 (n_37), .A2 (inputQ[5]), .A3 (inputQ[6]), .A4 (inputQ[7]));
INV_X1 i_65 (.ZN (n_33), .A (n_34));
NOR2_X1 i_64 (.ZN (n_32), .A1 (n_33), .A2 (inputQ[8]));
INV_X1 i_63 (.ZN (n_31), .A (n_32));
NOR2_X1 i_62 (.ZN (n_30), .A1 (n_31), .A2 (inputQ[9]));
NOR3_X1 i_61 (.ZN (n_29), .A1 (n_31), .A2 (inputQ[9]), .A3 (inputQ[10]));
INV_X1 i_60 (.ZN (n_28), .A (n_29));
NOR2_X1 i_59 (.ZN (n_27), .A1 (n_28), .A2 (inputQ[11]));
NOR3_X1 i_58 (.ZN (n_26), .A1 (n_28), .A2 (inputQ[11]), .A3 (inputQ[12]));
INV_X1 i_57 (.ZN (n_25), .A (n_26));
NOR2_X1 i_56 (.ZN (n_24), .A1 (n_25), .A2 (inputQ[13]));
NOR3_X1 i_55 (.ZN (n_23), .A1 (n_25), .A2 (inputQ[13]), .A3 (inputQ[14]));
INV_X1 i_54 (.ZN (n_22), .A (n_23));
NOR2_X1 i_53 (.ZN (n_21), .A1 (n_22), .A2 (inputQ[15]));
NOR3_X1 i_52 (.ZN (n_20), .A1 (n_22), .A2 (inputQ[15]), .A3 (inputQ[16]));
INV_X1 i_51 (.ZN (n_19), .A (n_20));
NOR2_X1 i_50 (.ZN (n_18), .A1 (n_19), .A2 (inputQ[17]));
NOR3_X1 i_49 (.ZN (n_17), .A1 (n_19), .A2 (inputQ[17]), .A3 (inputQ[18]));
INV_X1 i_48 (.ZN (n_16), .A (n_17));
NOR2_X1 i_47 (.ZN (n_15), .A1 (n_16), .A2 (inputQ[19]));
NOR3_X1 i_46 (.ZN (n_14), .A1 (n_16), .A2 (inputQ[19]), .A3 (inputQ[20]));
INV_X1 i_45 (.ZN (n_13), .A (n_14));
NOR2_X1 i_44 (.ZN (n_12), .A1 (n_13), .A2 (inputQ[21]));
NOR3_X1 i_43 (.ZN (n_11), .A1 (n_13), .A2 (inputQ[21]), .A3 (inputQ[22]));
INV_X1 i_42 (.ZN (n_10), .A (n_11));
NOR2_X1 i_41 (.ZN (n_9), .A1 (n_10), .A2 (inputQ[23]));
NOR3_X1 i_40 (.ZN (n_8), .A1 (n_10), .A2 (inputQ[23]), .A3 (inputQ[24]));
NAND2_X1 i_39 (.ZN (n_7), .A1 (n_8), .A2 (n_41));
NOR3_X1 i_38 (.ZN (n_6), .A1 (n_7), .A2 (inputQ[26]), .A3 (inputQ[27]));
NAND2_X1 i_37 (.ZN (n_5), .A1 (n_6), .A2 (n_42));
NOR2_X1 i_36 (.ZN (n_4), .A1 (n_5), .A2 (inputQ[29]));
NOR3_X1 i_35 (.ZN (n_3), .A1 (n_5), .A2 (inputQ[29]), .A3 (inputQ[30]));
XNOR2_X1 i_34 (.ZN (inputQ_inv22[31]), .A (inputQ[31]), .B (n_3));
XNOR2_X1 i_33 (.ZN (inputQ_inv22[30]), .A (inputQ[30]), .B (n_4));
XOR2_X1 i_32 (.Z (inputQ_inv22[29]), .A (inputQ[29]), .B (n_5));
XNOR2_X1 i_31 (.ZN (inputQ_inv22[28]), .A (inputQ[28]), .B (n_6));
OAI21_X1 i_30 (.ZN (n_2), .A (inputQ[27]), .B1 (n_7), .B2 (inputQ[26]));
INV_X1 i_29 (.ZN (n_1), .A (n_2));
NOR2_X1 i_28 (.ZN (inputQ_inv22[27]), .A1 (n_6), .A2 (n_1));
XOR2_X1 i_27 (.Z (inputQ_inv22[26]), .A (inputQ[26]), .B (n_7));
XNOR2_X1 i_26 (.ZN (inputQ_inv22[25]), .A (inputQ[25]), .B (n_8));
XNOR2_X1 i_25 (.ZN (inputQ_inv22[24]), .A (inputQ[24]), .B (n_9));
XNOR2_X1 i_24 (.ZN (inputQ_inv22[23]), .A (inputQ[23]), .B (n_11));
XNOR2_X1 i_23 (.ZN (inputQ_inv22[22]), .A (inputQ[22]), .B (n_12));
XNOR2_X1 i_22 (.ZN (inputQ_inv22[21]), .A (inputQ[21]), .B (n_14));
XNOR2_X1 i_21 (.ZN (inputQ_inv22[20]), .A (inputQ[20]), .B (n_15));
XNOR2_X1 i_20 (.ZN (inputQ_inv22[19]), .A (inputQ[19]), .B (n_17));
XNOR2_X1 i_19 (.ZN (inputQ_inv22[18]), .A (inputQ[18]), .B (n_18));
XNOR2_X1 i_18 (.ZN (inputQ_inv22[17]), .A (inputQ[17]), .B (n_20));
XNOR2_X1 i_17 (.ZN (inputQ_inv22[16]), .A (inputQ[16]), .B (n_21));
XNOR2_X1 i_16 (.ZN (inputQ_inv22[15]), .A (inputQ[15]), .B (n_23));
XNOR2_X1 i_15 (.ZN (inputQ_inv22[14]), .A (inputQ[14]), .B (n_24));
XNOR2_X1 i_14 (.ZN (inputQ_inv22[13]), .A (inputQ[13]), .B (n_26));
XNOR2_X1 i_13 (.ZN (inputQ_inv22[12]), .A (inputQ[12]), .B (n_27));
XNOR2_X1 i_12 (.ZN (inputQ_inv22[11]), .A (inputQ[11]), .B (n_29));
XNOR2_X1 i_11 (.ZN (inputQ_inv22[10]), .A (inputQ[10]), .B (n_30));
XNOR2_X1 i_10 (.ZN (inputQ_inv22[9]), .A (inputQ[9]), .B (n_32));
XNOR2_X1 i_9 (.ZN (inputQ_inv22[8]), .A (inputQ[8]), .B (n_34));
XNOR2_X1 i_8 (.ZN (inputQ_inv22[7]), .A (inputQ[7]), .B (n_35));
XNOR2_X1 i_7 (.ZN (inputQ_inv22[6]), .A (inputQ[6]), .B (n_36));
XOR2_X1 i_6 (.Z (inputQ_inv22[5]), .A (inputQ[5]), .B (n_37));
XOR2_X1 i_5 (.Z (inputQ_inv22[4]), .A (inputQ[4]), .B (n_38));
XOR2_X1 i_4 (.Z (inputQ_inv22[3]), .A (inputQ[3]), .B (n_39));
XOR2_X1 i_3 (.Z (inputQ_inv22[2]), .A (inputQ[2]), .B (n_40));
OAI21_X1 i_2 (.ZN (n_0), .A (inputQ[1]), .B1 (n_43), .B2 (inputQ[0]));
AND2_X1 i_1 (.ZN (inputQ_inv22[1]), .A1 (n_40), .A2 (n_0));
XNOR2_X1 i_0 (.ZN (inputQ_inv22[0]), .A (input_plus), .B (inputQ[0]));

endmodule //datapath__0_27

module registerNbits__parameterized0 (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [63:0] out;
input clk;
input en;
input [63:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_10;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire hfn_ipo_n5;
wire CTS_n_tid1_11;


AND2_X1 i_0_65 (.ZN (n_65), .A1 (hfn_ipo_n5), .A2 (inp[63]));
AND2_X1 i_0_64 (.ZN (n_64), .A1 (hfn_ipo_n5), .A2 (inp[62]));
AND2_X1 i_0_63 (.ZN (n_63), .A1 (hfn_ipo_n5), .A2 (inp[61]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (hfn_ipo_n5), .A2 (inp[60]));
AND2_X1 i_0_61 (.ZN (n_61), .A1 (hfn_ipo_n5), .A2 (inp[59]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (hfn_ipo_n5), .A2 (inp[58]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (hfn_ipo_n5), .A2 (inp[57]));
AND2_X1 i_0_58 (.ZN (n_58), .A1 (hfn_ipo_n5), .A2 (inp[56]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (hfn_ipo_n5), .A2 (inp[55]));
AND2_X1 i_0_56 (.ZN (n_56), .A1 (hfn_ipo_n5), .A2 (inp[54]));
AND2_X1 i_0_55 (.ZN (n_55), .A1 (hfn_ipo_n5), .A2 (inp[53]));
AND2_X1 i_0_54 (.ZN (n_54), .A1 (hfn_ipo_n5), .A2 (inp[52]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (hfn_ipo_n5), .A2 (inp[51]));
AND2_X1 i_0_52 (.ZN (n_52), .A1 (hfn_ipo_n5), .A2 (inp[50]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (hfn_ipo_n5), .A2 (inp[49]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (hfn_ipo_n5), .A2 (inp[48]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (hfn_ipo_n5), .A2 (inp[47]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (hfn_ipo_n5), .A2 (inp[46]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (hfn_ipo_n5), .A2 (inp[45]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (hfn_ipo_n5), .A2 (inp[44]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (hfn_ipo_n5), .A2 (inp[43]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (hfn_ipo_n5), .A2 (inp[42]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (hfn_ipo_n5), .A2 (inp[41]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (hfn_ipo_n5), .A2 (inp[40]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (hfn_ipo_n5), .A2 (inp[39]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (n_0_0), .A2 (inp[38]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (n_0_0), .A2 (inp[37]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (n_0_0), .A2 (inp[36]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (n_0_0), .A2 (inp[35]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (n_0_0), .A2 (inp[34]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (n_0_0), .A2 (inp[33]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (n_0_0), .A2 (inp[32]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (hfn_ipo_n5), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (hfn_ipo_n5), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (hfn_ipo_n5), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (hfn_ipo_n5), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (hfn_ipo_n5), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (hfn_ipo_n5), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (hfn_ipo_n5), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (hfn_ipo_n5), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (hfn_ipo_n5), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (hfn_ipo_n5), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (hfn_ipo_n5), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (hfn_ipo_n5), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (hfn_ipo_n5), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (hfn_ipo_n5), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (hfn_ipo_n5), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_10), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_10), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_10), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_10), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_10), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_10), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_10), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_10), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_10), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_10), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_10), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_10), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_10), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_10), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_10), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_10), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_10), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_10), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_10), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_10), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_10), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_10), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_10), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_10), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_10), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_10), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_10), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_10), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_10), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_10), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_10), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_10), .D (n_33));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n_tid1_10), .D (n_34));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n_tid1_10), .D (n_35));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n_tid1_10), .D (n_36));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n_tid1_10), .D (n_37));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n_tid1_10), .D (n_38));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n_tid1_10), .D (n_39));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n_tid1_10), .D (n_40));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n_tid1_10), .D (n_41));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n_tid1_10), .D (n_42));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n_tid1_10), .D (n_43));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n_tid1_10), .D (n_44));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n_tid1_10), .D (n_45));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n_tid1_10), .D (n_46));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n_tid1_10), .D (n_47));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n_tid1_10), .D (n_48));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n_tid1_10), .D (n_49));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n_tid1_10), .D (n_50));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n_tid1_10), .D (n_51));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n_tid1_10), .D (n_52));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n_tid1_10), .D (n_53));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n_tid1_10), .D (n_54));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n_tid1_10), .D (n_55));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n_tid1_10), .D (n_56));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n_tid1_10), .D (n_57));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n_tid1_10), .D (n_58));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n_tid1_10), .D (n_59));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n_tid1_10), .D (n_60));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n_tid1_10), .D (n_61));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n_tid1_10), .D (n_62));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n_tid1_10), .D (n_63));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (CTS_n_tid1_10), .D (n_64));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n_tid1_10), .D (n_65));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid1_11), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
BUF_X2 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_0_0));
CLKBUF_X3 CTS_L3_c_tid1_11 (.Z (CTS_n_tid1_10), .A (CTS_n_tid1_11));

endmodule //registerNbits__parameterized0

module datapath__0_17 (Acc, inputM_wire, p_0);

output [32:0] p_0;
input [31:0] Acc;
input [31:0] inputM_wire;
wire n_74;
wire n_100;
wire n_96;
wire n_0;
wire n_101;
wire n_97;
wire n_76;
wire n_72;
wire n_71;
wire n_69;
wire n_68;
wire n_66;
wire n_65;
wire n_63;
wire n_62;
wire n_60;
wire n_59;
wire n_57;
wire n_56;
wire n_54;
wire n_53;
wire n_51;
wire n_50;
wire n_48;
wire n_47;
wire n_45;
wire n_44;
wire n_42;
wire n_41;
wire n_39;
wire n_38;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_1;
wire n_102;
wire n_98;
wire n_79;
wire n_31;
wire n_30;
wire n_28;
wire n_27;
wire n_25;
wire n_24;
wire n_22;
wire n_21;
wire n_2;
wire n_81;
wire n_83;
wire n_20;
wire n_19;
wire n_3;
wire n_84;
wire n_85;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_4;
wire n_88;
wire n_90;
wire n_13;
wire n_12;
wire n_5;
wire n_92;
wire n_94;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_6;
wire n_103;
wire n_99;
wire n_7;
wire n_95;
wire n_93;
wire n_91;
wire n_89;
wire n_87;
wire n_86;
wire n_18;
wire n_82;
wire n_80;
wire n_23;
wire n_26;
wire n_29;
wire n_78;
wire n_32;
wire n_77;
wire n_37;
wire n_40;
wire n_43;
wire n_46;
wire n_49;
wire n_52;
wire n_55;
wire n_58;
wire n_61;
wire n_64;
wire n_67;
wire n_70;
wire n_75;
wire n_73;


INV_X1 i_136 (.ZN (n_103), .A (Acc[31]));
INV_X1 i_135 (.ZN (n_102), .A (Acc[16]));
INV_X1 i_134 (.ZN (n_101), .A (Acc[1]));
INV_X1 i_133 (.ZN (n_100), .A (Acc[0]));
INV_X1 i_132 (.ZN (n_99), .A (inputM_wire[31]));
INV_X1 i_131 (.ZN (n_98), .A (inputM_wire[16]));
INV_X1 i_130 (.ZN (n_97), .A (inputM_wire[1]));
INV_X1 i_129 (.ZN (n_96), .A (inputM_wire[0]));
NAND2_X1 i_128 (.ZN (n_95), .A1 (Acc[30]), .A2 (inputM_wire[30]));
XNOR2_X1 i_127 (.ZN (n_94), .A (Acc[29]), .B (inputM_wire[29]));
INV_X1 i_126 (.ZN (n_93), .A (n_94));
NAND2_X1 i_125 (.ZN (n_92), .A1 (Acc[28]), .A2 (inputM_wire[28]));
NOR2_X1 i_124 (.ZN (n_91), .A1 (Acc[28]), .A2 (inputM_wire[28]));
XNOR2_X1 i_123 (.ZN (n_90), .A (Acc[27]), .B (inputM_wire[27]));
INV_X1 i_122 (.ZN (n_89), .A (n_90));
NAND2_X1 i_121 (.ZN (n_88), .A1 (Acc[26]), .A2 (inputM_wire[26]));
NOR2_X1 i_120 (.ZN (n_87), .A1 (Acc[26]), .A2 (inputM_wire[26]));
NAND2_X1 i_119 (.ZN (n_86), .A1 (Acc[24]), .A2 (inputM_wire[24]));
OAI21_X1 i_118 (.ZN (n_85), .A (n_86), .B1 (Acc[24]), .B2 (inputM_wire[24]));
NAND2_X1 i_117 (.ZN (n_84), .A1 (Acc[23]), .A2 (inputM_wire[23]));
XNOR2_X1 i_116 (.ZN (n_83), .A (Acc[22]), .B (inputM_wire[22]));
INV_X1 i_115 (.ZN (n_82), .A (n_83));
NAND2_X1 i_114 (.ZN (n_81), .A1 (Acc[21]), .A2 (inputM_wire[21]));
NOR2_X1 i_113 (.ZN (n_80), .A1 (Acc[21]), .A2 (inputM_wire[21]));
XNOR2_X1 i_112 (.ZN (n_79), .A (Acc[17]), .B (inputM_wire[17]));
INV_X1 i_111 (.ZN (n_78), .A (n_79));
NAND2_X1 i_110 (.ZN (n_77), .A1 (Acc[15]), .A2 (inputM_wire[15]));
XNOR2_X1 i_109 (.ZN (n_76), .A (Acc[2]), .B (inputM_wire[2]));
INV_X1 i_108 (.ZN (n_75), .A (n_76));
NOR2_X1 i_107 (.ZN (n_74), .A1 (n_100), .A2 (n_96));
AOI21_X1 i_106 (.ZN (n_73), .A (n_74), .B1 (Acc[1]), .B2 (inputM_wire[1]));
AOI21_X1 i_105 (.ZN (n_72), .A (n_73), .B1 (n_101), .B2 (n_97));
AOI22_X1 i_104 (.ZN (n_71), .A1 (Acc[2]), .A2 (inputM_wire[2]), .B1 (n_75), .B2 (n_72));
INV_X1 i_103 (.ZN (n_70), .A (n_71));
XOR2_X1 i_102 (.Z (n_69), .A (Acc[3]), .B (inputM_wire[3]));
AOI22_X1 i_101 (.ZN (n_68), .A1 (Acc[3]), .A2 (inputM_wire[3]), .B1 (n_70), .B2 (n_69));
INV_X1 i_100 (.ZN (n_67), .A (n_68));
XOR2_X1 i_99 (.Z (n_66), .A (Acc[4]), .B (inputM_wire[4]));
AOI22_X1 i_98 (.ZN (n_65), .A1 (Acc[4]), .A2 (inputM_wire[4]), .B1 (n_67), .B2 (n_66));
INV_X1 i_97 (.ZN (n_64), .A (n_65));
XOR2_X1 i_96 (.Z (n_63), .A (Acc[5]), .B (inputM_wire[5]));
AOI22_X1 i_95 (.ZN (n_62), .A1 (Acc[5]), .A2 (inputM_wire[5]), .B1 (n_64), .B2 (n_63));
INV_X1 i_94 (.ZN (n_61), .A (n_62));
XOR2_X1 i_93 (.Z (n_60), .A (Acc[6]), .B (inputM_wire[6]));
AOI22_X1 i_92 (.ZN (n_59), .A1 (Acc[6]), .A2 (inputM_wire[6]), .B1 (n_61), .B2 (n_60));
INV_X1 i_91 (.ZN (n_58), .A (n_59));
XOR2_X1 i_90 (.Z (n_57), .A (Acc[7]), .B (inputM_wire[7]));
AOI22_X1 i_89 (.ZN (n_56), .A1 (Acc[7]), .A2 (inputM_wire[7]), .B1 (n_58), .B2 (n_57));
INV_X1 i_88 (.ZN (n_55), .A (n_56));
XOR2_X1 i_87 (.Z (n_54), .A (Acc[8]), .B (inputM_wire[8]));
AOI22_X1 i_86 (.ZN (n_53), .A1 (Acc[8]), .A2 (inputM_wire[8]), .B1 (n_55), .B2 (n_54));
INV_X1 i_85 (.ZN (n_52), .A (n_53));
XOR2_X1 i_84 (.Z (n_51), .A (Acc[9]), .B (inputM_wire[9]));
AOI22_X1 i_83 (.ZN (n_50), .A1 (Acc[9]), .A2 (inputM_wire[9]), .B1 (n_52), .B2 (n_51));
INV_X1 i_82 (.ZN (n_49), .A (n_50));
XOR2_X1 i_81 (.Z (n_48), .A (Acc[10]), .B (inputM_wire[10]));
AOI22_X1 i_80 (.ZN (n_47), .A1 (Acc[10]), .A2 (inputM_wire[10]), .B1 (n_49), .B2 (n_48));
INV_X1 i_79 (.ZN (n_46), .A (n_47));
XOR2_X1 i_78 (.Z (n_45), .A (Acc[11]), .B (inputM_wire[11]));
AOI22_X1 i_77 (.ZN (n_44), .A1 (Acc[11]), .A2 (inputM_wire[11]), .B1 (n_46), .B2 (n_45));
INV_X1 i_76 (.ZN (n_43), .A (n_44));
XOR2_X1 i_75 (.Z (n_42), .A (Acc[12]), .B (inputM_wire[12]));
AOI22_X1 i_74 (.ZN (n_41), .A1 (Acc[12]), .A2 (inputM_wire[12]), .B1 (n_43), .B2 (n_42));
INV_X1 i_73 (.ZN (n_40), .A (n_41));
XOR2_X1 i_72 (.Z (n_39), .A (Acc[13]), .B (inputM_wire[13]));
AOI22_X1 i_71 (.ZN (n_38), .A1 (Acc[13]), .A2 (inputM_wire[13]), .B1 (n_40), .B2 (n_39));
INV_X1 i_70 (.ZN (n_37), .A (n_38));
XOR2_X1 i_69 (.Z (n_36), .A (Acc[14]), .B (inputM_wire[14]));
AOI22_X1 i_68 (.ZN (n_35), .A1 (Acc[14]), .A2 (inputM_wire[14]), .B1 (n_37), .B2 (n_36));
OAI21_X1 i_67 (.ZN (n_34), .A (n_77), .B1 (Acc[15]), .B2 (inputM_wire[15]));
OAI21_X1 i_66 (.ZN (n_33), .A (n_77), .B1 (n_35), .B2 (n_34));
OAI21_X1 i_65 (.ZN (n_32), .A (n_33), .B1 (Acc[16]), .B2 (inputM_wire[16]));
OAI21_X1 i_64 (.ZN (n_31), .A (n_32), .B1 (n_102), .B2 (n_98));
AOI22_X1 i_63 (.ZN (n_30), .A1 (Acc[17]), .A2 (inputM_wire[17]), .B1 (n_78), .B2 (n_31));
INV_X1 i_62 (.ZN (n_29), .A (n_30));
XOR2_X1 i_61 (.Z (n_28), .A (Acc[18]), .B (inputM_wire[18]));
AOI22_X1 i_60 (.ZN (n_27), .A1 (Acc[18]), .A2 (inputM_wire[18]), .B1 (n_29), .B2 (n_28));
INV_X1 i_59 (.ZN (n_26), .A (n_27));
XOR2_X1 i_58 (.Z (n_25), .A (Acc[19]), .B (inputM_wire[19]));
AOI22_X1 i_57 (.ZN (n_24), .A1 (Acc[19]), .A2 (inputM_wire[19]), .B1 (n_26), .B2 (n_25));
INV_X1 i_56 (.ZN (n_23), .A (n_24));
XOR2_X1 i_55 (.Z (n_22), .A (Acc[20]), .B (inputM_wire[20]));
AOI22_X1 i_54 (.ZN (n_21), .A1 (Acc[20]), .A2 (inputM_wire[20]), .B1 (n_23), .B2 (n_22));
AOI21_X1 i_53 (.ZN (n_20), .A (n_80), .B1 (n_81), .B2 (n_21));
AOI22_X1 i_52 (.ZN (n_19), .A1 (Acc[22]), .A2 (inputM_wire[22]), .B1 (n_82), .B2 (n_20));
NAND2_X1 i_51 (.ZN (n_18), .A1 (n_84), .A2 (n_19));
OAI21_X1 i_50 (.ZN (n_17), .A (n_18), .B1 (Acc[23]), .B2 (inputM_wire[23]));
OAI21_X1 i_49 (.ZN (n_16), .A (n_86), .B1 (n_85), .B2 (n_17));
XOR2_X1 i_48 (.Z (n_15), .A (Acc[25]), .B (inputM_wire[25]));
AOI22_X1 i_47 (.ZN (n_14), .A1 (Acc[25]), .A2 (inputM_wire[25]), .B1 (n_16), .B2 (n_15));
AOI21_X1 i_46 (.ZN (n_13), .A (n_87), .B1 (n_88), .B2 (n_14));
AOI22_X1 i_45 (.ZN (n_12), .A1 (Acc[27]), .A2 (inputM_wire[27]), .B1 (n_89), .B2 (n_13));
AOI21_X1 i_44 (.ZN (n_11), .A (n_91), .B1 (n_92), .B2 (n_12));
AOI22_X1 i_43 (.ZN (n_10), .A1 (Acc[29]), .A2 (inputM_wire[29]), .B1 (n_93), .B2 (n_11));
OAI21_X1 i_42 (.ZN (n_9), .A (n_95), .B1 (Acc[30]), .B2 (inputM_wire[30]));
OAI21_X1 i_41 (.ZN (n_8), .A (n_95), .B1 (n_10), .B2 (n_9));
AOI21_X1 i_40 (.ZN (n_7), .A (n_8), .B1 (Acc[31]), .B2 (inputM_wire[31]));
AOI21_X1 i_39 (.ZN (p_0[32]), .A (n_7), .B1 (n_103), .B2 (n_99));
OAI22_X1 i_38 (.ZN (n_6), .A1 (n_103), .A2 (n_99), .B1 (Acc[31]), .B2 (inputM_wire[31]));
XNOR2_X1 i_37 (.ZN (p_0[31]), .A (n_8), .B (n_6));
XOR2_X1 i_36 (.Z (p_0[30]), .A (n_10), .B (n_9));
XNOR2_X1 i_35 (.ZN (p_0[29]), .A (n_94), .B (n_11));
OAI21_X1 i_34 (.ZN (n_5), .A (n_92), .B1 (Acc[28]), .B2 (inputM_wire[28]));
XOR2_X1 i_33 (.Z (p_0[28]), .A (n_12), .B (n_5));
XNOR2_X1 i_32 (.ZN (p_0[27]), .A (n_90), .B (n_13));
OAI21_X1 i_31 (.ZN (n_4), .A (n_88), .B1 (Acc[26]), .B2 (inputM_wire[26]));
XOR2_X1 i_30 (.Z (p_0[26]), .A (n_14), .B (n_4));
XOR2_X1 i_29 (.Z (p_0[25]), .A (n_16), .B (n_15));
XOR2_X1 i_28 (.Z (p_0[24]), .A (n_85), .B (n_17));
OAI21_X1 i_27 (.ZN (n_3), .A (n_84), .B1 (Acc[23]), .B2 (inputM_wire[23]));
XOR2_X1 i_26 (.Z (p_0[23]), .A (n_19), .B (n_3));
XNOR2_X1 i_25 (.ZN (p_0[22]), .A (n_83), .B (n_20));
OAI21_X1 i_24 (.ZN (n_2), .A (n_81), .B1 (Acc[21]), .B2 (inputM_wire[21]));
XOR2_X1 i_23 (.Z (p_0[21]), .A (n_21), .B (n_2));
XNOR2_X1 i_22 (.ZN (p_0[20]), .A (n_24), .B (n_22));
XNOR2_X1 i_21 (.ZN (p_0[19]), .A (n_27), .B (n_25));
XNOR2_X1 i_20 (.ZN (p_0[18]), .A (n_30), .B (n_28));
XNOR2_X1 i_19 (.ZN (p_0[17]), .A (n_79), .B (n_31));
OAI22_X1 i_18 (.ZN (n_1), .A1 (Acc[16]), .A2 (inputM_wire[16]), .B1 (n_102), .B2 (n_98));
XNOR2_X1 i_17 (.ZN (p_0[16]), .A (n_33), .B (n_1));
XOR2_X1 i_16 (.Z (p_0[15]), .A (n_35), .B (n_34));
XNOR2_X1 i_15 (.ZN (p_0[14]), .A (n_38), .B (n_36));
XNOR2_X1 i_14 (.ZN (p_0[13]), .A (n_41), .B (n_39));
XNOR2_X1 i_13 (.ZN (p_0[12]), .A (n_44), .B (n_42));
XNOR2_X1 i_12 (.ZN (p_0[11]), .A (n_47), .B (n_45));
XNOR2_X1 i_11 (.ZN (p_0[10]), .A (n_50), .B (n_48));
XNOR2_X1 i_10 (.ZN (p_0[9]), .A (n_53), .B (n_51));
XNOR2_X1 i_9 (.ZN (p_0[8]), .A (n_56), .B (n_54));
XNOR2_X1 i_8 (.ZN (p_0[7]), .A (n_59), .B (n_57));
XNOR2_X1 i_7 (.ZN (p_0[6]), .A (n_62), .B (n_60));
XNOR2_X1 i_6 (.ZN (p_0[5]), .A (n_65), .B (n_63));
XNOR2_X1 i_5 (.ZN (p_0[4]), .A (n_68), .B (n_66));
XNOR2_X1 i_4 (.ZN (p_0[3]), .A (n_71), .B (n_69));
XNOR2_X1 i_3 (.ZN (p_0[2]), .A (n_76), .B (n_72));
OAI22_X1 i_2 (.ZN (n_0), .A1 (n_101), .A2 (n_97), .B1 (Acc[1]), .B2 (inputM_wire[1]));
XNOR2_X1 i_1 (.ZN (p_0[1]), .A (n_74), .B (n_0));
AOI21_X1 i_0 (.ZN (p_0[0]), .A (n_74), .B1 (n_100), .B2 (n_96));

endmodule //datapath__0_17

module datapath (input_plus, p_0, p_1);

output [63:0] p_0;
input input_plus;
input [63:0] p_1;
wire CLOCK_slh_n5;
wire n_86;
wire n_0;
wire n_92;
wire n_85;
wire n_84;
wire n_83;
wire n_81;
wire n_1;
wire n_82;
wire n_80;
wire n_2;
wire n_88;
wire n_87;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_74;
wire n_73;
wire n_71;
wire n_70;
wire n_68;
wire n_67;
wire n_65;
wire n_64;
wire n_62;
wire n_61;
wire n_59;
wire n_58;
wire n_56;
wire n_55;
wire n_53;
wire n_52;
wire n_50;
wire n_49;
wire n_47;
wire n_46;
wire n_44;
wire n_43;
wire n_41;
wire n_40;
wire n_38;
wire n_37;
wire n_35;
wire n_34;
wire n_32;
wire n_31;
wire n_29;
wire n_28;
wire n_26;
wire n_25;
wire n_23;
wire n_22;
wire n_20;
wire n_19;
wire n_17;
wire n_16;
wire n_14;
wire n_13;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_3;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_91;
wire n_90;
wire n_12;
wire n_15;
wire n_18;
wire n_21;
wire n_24;
wire n_27;
wire n_30;
wire n_33;
wire n_36;
wire n_39;
wire n_42;
wire n_45;
wire n_48;
wire n_51;
wire n_54;
wire n_57;
wire n_60;
wire n_63;
wire n_66;
wire n_69;
wire n_72;
wire n_75;
wire n_89;


INV_X1 i_156 (.ZN (n_92), .A (CLOCK_slh_n5));
INV_X1 i_155 (.ZN (n_91), .A (p_1[60]));
INV_X1 i_154 (.ZN (n_90), .A (p_1[57]));
INV_X1 i_153 (.ZN (n_89), .A (p_1[9]));
INV_X1 i_152 (.ZN (n_88), .A (p_1[8]));
INV_X1 i_151 (.ZN (n_87), .A (p_1[7]));
OR3_X1 i_150 (.ZN (n_86), .A1 (n_92), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_149 (.ZN (n_85), .A1 (n_86), .A2 (p_1[2]));
OR2_X1 i_148 (.ZN (n_84), .A1 (n_85), .A2 (p_1[3]));
OR2_X1 i_147 (.ZN (n_83), .A1 (n_84), .A2 (p_1[4]));
NOR3_X1 i_146 (.ZN (n_82), .A1 (n_83), .A2 (p_1[5]), .A3 (p_1[6]));
INV_X1 i_145 (.ZN (n_81), .A (n_82));
NOR3_X1 i_144 (.ZN (n_80), .A1 (n_81), .A2 (p_1[7]), .A3 (p_1[8]));
NAND2_X1 i_143 (.ZN (n_79), .A1 (n_80), .A2 (n_89));
NOR2_X1 i_142 (.ZN (n_78), .A1 (n_79), .A2 (p_1[10]));
NOR3_X1 i_141 (.ZN (n_77), .A1 (n_79), .A2 (p_1[10]), .A3 (p_1[11]));
NOR4_X1 i_140 (.ZN (n_76), .A1 (n_79), .A2 (p_1[10]), .A3 (p_1[11]), .A4 (p_1[12]));
INV_X1 i_139 (.ZN (n_75), .A (n_76));
NOR2_X1 i_138 (.ZN (n_74), .A1 (n_75), .A2 (p_1[13]));
NOR3_X1 i_137 (.ZN (n_73), .A1 (n_75), .A2 (p_1[13]), .A3 (p_1[14]));
INV_X1 i_136 (.ZN (n_72), .A (n_73));
NOR2_X1 i_135 (.ZN (n_71), .A1 (n_72), .A2 (p_1[15]));
NOR3_X1 i_134 (.ZN (n_70), .A1 (n_72), .A2 (p_1[15]), .A3 (p_1[16]));
INV_X1 i_133 (.ZN (n_69), .A (n_70));
NOR2_X1 i_132 (.ZN (n_68), .A1 (n_69), .A2 (p_1[17]));
NOR3_X1 i_131 (.ZN (n_67), .A1 (n_69), .A2 (p_1[17]), .A3 (p_1[18]));
INV_X1 i_130 (.ZN (n_66), .A (n_67));
NOR2_X1 i_129 (.ZN (n_65), .A1 (n_66), .A2 (p_1[19]));
NOR3_X1 i_128 (.ZN (n_64), .A1 (n_66), .A2 (p_1[19]), .A3 (p_1[20]));
INV_X1 i_127 (.ZN (n_63), .A (n_64));
NOR2_X1 i_126 (.ZN (n_62), .A1 (n_63), .A2 (p_1[21]));
NOR3_X1 i_125 (.ZN (n_61), .A1 (n_63), .A2 (p_1[21]), .A3 (p_1[22]));
INV_X1 i_124 (.ZN (n_60), .A (n_61));
NOR2_X1 i_123 (.ZN (n_59), .A1 (n_60), .A2 (p_1[23]));
NOR3_X1 i_122 (.ZN (n_58), .A1 (n_60), .A2 (p_1[23]), .A3 (p_1[24]));
INV_X1 i_121 (.ZN (n_57), .A (n_58));
NOR2_X1 i_120 (.ZN (n_56), .A1 (n_57), .A2 (p_1[25]));
NOR3_X1 i_119 (.ZN (n_55), .A1 (n_57), .A2 (p_1[25]), .A3 (p_1[26]));
INV_X1 i_118 (.ZN (n_54), .A (n_55));
NOR2_X1 i_117 (.ZN (n_53), .A1 (n_54), .A2 (p_1[27]));
NOR3_X1 i_116 (.ZN (n_52), .A1 (n_54), .A2 (p_1[27]), .A3 (p_1[28]));
INV_X1 i_115 (.ZN (n_51), .A (n_52));
NOR2_X1 i_114 (.ZN (n_50), .A1 (n_51), .A2 (p_1[29]));
NOR3_X1 i_113 (.ZN (n_49), .A1 (n_51), .A2 (p_1[29]), .A3 (p_1[30]));
INV_X1 i_112 (.ZN (n_48), .A (n_49));
NOR2_X1 i_111 (.ZN (n_47), .A1 (n_48), .A2 (p_1[31]));
NOR3_X1 i_110 (.ZN (n_46), .A1 (n_48), .A2 (p_1[31]), .A3 (p_1[32]));
INV_X1 i_109 (.ZN (n_45), .A (n_46));
NOR2_X1 i_108 (.ZN (n_44), .A1 (n_45), .A2 (p_1[33]));
NOR3_X1 i_107 (.ZN (n_43), .A1 (n_45), .A2 (p_1[33]), .A3 (p_1[34]));
INV_X1 i_106 (.ZN (n_42), .A (n_43));
NOR2_X1 i_105 (.ZN (n_41), .A1 (n_42), .A2 (p_1[35]));
NOR3_X1 i_104 (.ZN (n_40), .A1 (n_42), .A2 (p_1[35]), .A3 (p_1[36]));
INV_X1 i_103 (.ZN (n_39), .A (n_40));
NOR2_X1 i_102 (.ZN (n_38), .A1 (n_39), .A2 (p_1[37]));
NOR3_X1 i_101 (.ZN (n_37), .A1 (n_39), .A2 (p_1[37]), .A3 (p_1[38]));
INV_X1 i_100 (.ZN (n_36), .A (n_37));
NOR2_X1 i_99 (.ZN (n_35), .A1 (n_36), .A2 (p_1[39]));
NOR3_X1 i_98 (.ZN (n_34), .A1 (n_36), .A2 (p_1[39]), .A3 (p_1[40]));
INV_X1 i_97 (.ZN (n_33), .A (n_34));
NOR2_X1 i_96 (.ZN (n_32), .A1 (n_33), .A2 (p_1[41]));
NOR3_X1 i_95 (.ZN (n_31), .A1 (n_33), .A2 (p_1[41]), .A3 (p_1[42]));
INV_X1 i_94 (.ZN (n_30), .A (n_31));
NOR2_X1 i_93 (.ZN (n_29), .A1 (n_30), .A2 (p_1[43]));
NOR3_X1 i_92 (.ZN (n_28), .A1 (n_30), .A2 (p_1[43]), .A3 (p_1[44]));
INV_X1 i_91 (.ZN (n_27), .A (n_28));
NOR2_X1 i_90 (.ZN (n_26), .A1 (n_27), .A2 (p_1[45]));
NOR3_X1 i_89 (.ZN (n_25), .A1 (n_27), .A2 (p_1[45]), .A3 (p_1[46]));
INV_X1 i_88 (.ZN (n_24), .A (n_25));
NOR2_X1 i_87 (.ZN (n_23), .A1 (n_24), .A2 (p_1[47]));
NOR3_X1 i_86 (.ZN (n_22), .A1 (n_24), .A2 (p_1[47]), .A3 (p_1[48]));
INV_X1 i_85 (.ZN (n_21), .A (n_22));
NOR2_X1 i_84 (.ZN (n_20), .A1 (n_21), .A2 (p_1[49]));
NOR3_X1 i_83 (.ZN (n_19), .A1 (n_21), .A2 (p_1[49]), .A3 (p_1[50]));
INV_X1 i_82 (.ZN (n_18), .A (n_19));
NOR2_X1 i_81 (.ZN (n_17), .A1 (n_18), .A2 (p_1[51]));
NOR3_X1 i_80 (.ZN (n_16), .A1 (n_18), .A2 (p_1[51]), .A3 (p_1[52]));
INV_X1 i_79 (.ZN (n_15), .A (n_16));
NOR2_X1 i_78 (.ZN (n_14), .A1 (n_15), .A2 (p_1[53]));
NOR3_X1 i_77 (.ZN (n_13), .A1 (n_15), .A2 (p_1[53]), .A3 (p_1[54]));
INV_X1 i_76 (.ZN (n_12), .A (n_13));
NOR2_X1 i_75 (.ZN (n_11), .A1 (n_12), .A2 (p_1[55]));
NOR3_X1 i_74 (.ZN (n_10), .A1 (n_12), .A2 (p_1[55]), .A3 (p_1[56]));
NAND2_X1 i_73 (.ZN (n_9), .A1 (n_10), .A2 (n_90));
NOR3_X1 i_72 (.ZN (n_8), .A1 (n_9), .A2 (p_1[58]), .A3 (p_1[59]));
NAND2_X1 i_71 (.ZN (n_7), .A1 (n_8), .A2 (n_91));
NOR2_X1 i_70 (.ZN (n_6), .A1 (n_7), .A2 (p_1[61]));
NOR3_X1 i_69 (.ZN (n_5), .A1 (n_7), .A2 (p_1[61]), .A3 (p_1[62]));
XNOR2_X1 i_68 (.ZN (p_0[63]), .A (p_1[63]), .B (n_5));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (p_1[62]), .B (n_6));
XOR2_X1 i_66 (.Z (p_0[61]), .A (p_1[61]), .B (n_7));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (p_1[60]), .B (n_8));
OAI21_X1 i_64 (.ZN (n_4), .A (p_1[59]), .B1 (n_9), .B2 (p_1[58]));
INV_X1 i_63 (.ZN (n_3), .A (n_4));
NOR2_X1 i_62 (.ZN (p_0[59]), .A1 (n_8), .A2 (n_3));
XOR2_X1 i_61 (.Z (p_0[58]), .A (p_1[58]), .B (n_9));
XNOR2_X1 i_60 (.ZN (p_0[57]), .A (p_1[57]), .B (n_10));
XNOR2_X1 i_59 (.ZN (p_0[56]), .A (p_1[56]), .B (n_11));
XNOR2_X1 i_58 (.ZN (p_0[55]), .A (p_1[55]), .B (n_13));
XNOR2_X1 i_57 (.ZN (p_0[54]), .A (p_1[54]), .B (n_14));
XNOR2_X1 i_56 (.ZN (p_0[53]), .A (p_1[53]), .B (n_16));
XNOR2_X1 i_55 (.ZN (p_0[52]), .A (p_1[52]), .B (n_17));
XNOR2_X1 i_54 (.ZN (p_0[51]), .A (p_1[51]), .B (n_19));
XNOR2_X1 i_53 (.ZN (p_0[50]), .A (p_1[50]), .B (n_20));
XNOR2_X1 i_52 (.ZN (p_0[49]), .A (p_1[49]), .B (n_22));
XNOR2_X1 i_51 (.ZN (p_0[48]), .A (p_1[48]), .B (n_23));
XNOR2_X1 i_50 (.ZN (p_0[47]), .A (p_1[47]), .B (n_25));
XNOR2_X1 i_49 (.ZN (p_0[46]), .A (p_1[46]), .B (n_26));
XNOR2_X1 i_48 (.ZN (p_0[45]), .A (p_1[45]), .B (n_28));
XNOR2_X1 i_47 (.ZN (p_0[44]), .A (p_1[44]), .B (n_29));
XNOR2_X1 i_46 (.ZN (p_0[43]), .A (p_1[43]), .B (n_31));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (p_1[42]), .B (n_32));
XNOR2_X1 i_44 (.ZN (p_0[41]), .A (p_1[41]), .B (n_34));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (p_1[40]), .B (n_35));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (p_1[39]), .B (n_37));
XNOR2_X1 i_41 (.ZN (p_0[38]), .A (p_1[38]), .B (n_38));
XNOR2_X1 i_40 (.ZN (p_0[37]), .A (p_1[37]), .B (n_40));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (p_1[36]), .B (n_41));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (p_1[35]), .B (n_43));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (p_1[34]), .B (n_44));
XNOR2_X1 i_36 (.ZN (p_0[33]), .A (p_1[33]), .B (n_46));
XNOR2_X1 i_35 (.ZN (p_0[32]), .A (p_1[32]), .B (n_47));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (p_1[31]), .B (n_49));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (p_1[30]), .B (n_50));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (p_1[29]), .B (n_52));
XNOR2_X1 i_31 (.ZN (p_0[28]), .A (p_1[28]), .B (n_53));
XNOR2_X1 i_30 (.ZN (p_0[27]), .A (p_1[27]), .B (n_55));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (p_1[26]), .B (n_56));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_58));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_59));
XNOR2_X1 i_26 (.ZN (p_0[23]), .A (p_1[23]), .B (n_61));
XNOR2_X1 i_25 (.ZN (p_0[22]), .A (p_1[22]), .B (n_62));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_64));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_65));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_67));
XNOR2_X1 i_21 (.ZN (p_0[18]), .A (p_1[18]), .B (n_68));
XNOR2_X1 i_20 (.ZN (p_0[17]), .A (p_1[17]), .B (n_70));
XNOR2_X1 i_19 (.ZN (p_0[16]), .A (p_1[16]), .B (n_71));
XNOR2_X1 i_18 (.ZN (p_0[15]), .A (p_1[15]), .B (n_73));
XNOR2_X1 i_17 (.ZN (p_0[14]), .A (p_1[14]), .B (n_74));
XNOR2_X1 i_16 (.ZN (p_0[13]), .A (p_1[13]), .B (n_76));
XNOR2_X1 i_15 (.ZN (p_0[12]), .A (p_1[12]), .B (n_77));
XNOR2_X1 i_14 (.ZN (p_0[11]), .A (p_1[11]), .B (n_78));
XOR2_X1 i_13 (.Z (p_0[10]), .A (p_1[10]), .B (n_79));
XNOR2_X1 i_12 (.ZN (p_0[9]), .A (p_1[9]), .B (n_80));
AOI21_X1 i_11 (.ZN (n_2), .A (n_88), .B1 (n_82), .B2 (n_87));
NOR2_X1 i_10 (.ZN (p_0[8]), .A1 (n_80), .A2 (n_2));
XNOR2_X1 i_9 (.ZN (p_0[7]), .A (p_1[7]), .B (n_82));
OAI21_X1 i_8 (.ZN (n_1), .A (p_1[6]), .B1 (n_83), .B2 (p_1[5]));
AND2_X1 i_7 (.ZN (p_0[6]), .A1 (n_81), .A2 (n_1));
XOR2_X1 i_6 (.Z (p_0[5]), .A (p_1[5]), .B (n_83));
XOR2_X1 i_5 (.Z (p_0[4]), .A (p_1[4]), .B (n_84));
XOR2_X1 i_4 (.Z (p_0[3]), .A (p_1[3]), .B (n_85));
XOR2_X1 i_3 (.Z (p_0[2]), .A (p_1[2]), .B (n_86));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[1]), .B1 (n_92), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[1]), .A1 (n_86), .A2 (n_0));
XNOR2_X1 i_0 (.ZN (p_0[0]), .A (CLOCK_slh_n5), .B (p_1[0]));
CLKBUF_X1 CLOCK_slh__c1 (.Z (CLOCK_slh_n5), .A (input_plus));

endmodule //datapath

module controller (clk_CTS_0_PP_0, clk_CTS_0_PP_1, clk, reset, inputQ_wire, inputM_wire, 
    Mbit, Qbit, input_plus, out);

output [63:0] out;
output clk_CTS_0_PP_0;
input Mbit;
input Qbit;
input clk;
input [31:0] inputM_wire;
input [31:0] inputQ_wire;
input input_plus;
input reset;
input clk_CTS_0_PP_1;
wire CTS_n_tid0_198;
wire \inputQ_reg[31] ;
wire \inputQ_reg[30] ;
wire \inputQ_reg[29] ;
wire \inputQ_reg[28] ;
wire \inputQ_reg[27] ;
wire \inputQ_reg[26] ;
wire \inputQ_reg[25] ;
wire \inputQ_reg[24] ;
wire \inputQ_reg[23] ;
wire \inputQ_reg[22] ;
wire \inputQ_reg[21] ;
wire \inputQ_reg[20] ;
wire \inputQ_reg[19] ;
wire \inputQ_reg[18] ;
wire \inputQ_reg[17] ;
wire \inputQ_reg[16] ;
wire \inputQ_reg[15] ;
wire \inputQ_reg[14] ;
wire \inputQ_reg[13] ;
wire \inputQ_reg[12] ;
wire \inputQ_reg[11] ;
wire \inputQ_reg[10] ;
wire \inputQ_reg[9] ;
wire \inputQ_reg[8] ;
wire \inputQ_reg[7] ;
wire \inputQ_reg[6] ;
wire \inputQ_reg[5] ;
wire \inputQ_reg[4] ;
wire \inputQ_reg[3] ;
wire \inputQ_reg[2] ;
wire \inputQ_reg[1] ;
wire \inputQ_reg[0] ;
wire \Acc[31] ;
wire \Acc[30] ;
wire \Acc[29] ;
wire \Acc[28] ;
wire \Acc[27] ;
wire \Acc[26] ;
wire \Acc[25] ;
wire \Acc[24] ;
wire \Acc[23] ;
wire \Acc[22] ;
wire \Acc[21] ;
wire \Acc[20] ;
wire \Acc[19] ;
wire \Acc[18] ;
wire \Acc[17] ;
wire \Acc[16] ;
wire \Acc[15] ;
wire \Acc[14] ;
wire \Acc[13] ;
wire \Acc[12] ;
wire \Acc[11] ;
wire \Acc[10] ;
wire \Acc[9] ;
wire \Acc[8] ;
wire \Acc[7] ;
wire \Acc[6] ;
wire \Acc[5] ;
wire \Acc[4] ;
wire \Acc[3] ;
wire \Acc[2] ;
wire \Acc[1] ;
wire \Acc[0] ;
wire CTS_n_tid0_121;
wire CTS_n_tid0_209;
wire CTS_n_tid0_188;
wire CTS_n_tid0_49;
wire CTS_n_tid0_56;
wire CTS_n_tid0_122;
wire CTS_n_tid1_17;
wire hfn_ipo_n12;
wire hfn_ipo_n11;
wire hfn_ipo_n10;
wire hfn_ipo_n9;
wire \count[5] ;
wire \count[4] ;
wire \count[3] ;
wire \count[2] ;
wire \count[1] ;
wire \count[0] ;
wire \state[2] ;
wire \state[1] ;
wire \state[0] ;
wire \add_output[31] ;
wire \add_output[30] ;
wire \add_output[29] ;
wire \add_output[28] ;
wire \add_output[27] ;
wire \add_output[26] ;
wire \add_output[25] ;
wire \add_output[24] ;
wire \add_output[23] ;
wire \add_output[22] ;
wire \add_output[21] ;
wire \add_output[20] ;
wire \add_output[19] ;
wire \add_output[18] ;
wire \add_output[17] ;
wire \add_output[16] ;
wire \add_output[15] ;
wire \add_output[14] ;
wire \add_output[13] ;
wire \add_output[12] ;
wire \add_output[11] ;
wire \add_output[10] ;
wire \add_output[9] ;
wire \add_output[8] ;
wire \add_output[7] ;
wire \add_output[6] ;
wire \add_output[5] ;
wire \add_output[4] ;
wire \add_output[3] ;
wire \add_output[2] ;
wire \add_output[1] ;
wire \add_output[0] ;
wire lsb_reg;
wire c_output;
wire start;
wire n_2_0;
wire n_2_1;
wire n_2_2;
wire n_2_3;
wire n_2_4;
wire n_2_5;
wire n_2_6;
wire n_2_7;
wire n_2_8;
wire n_2_9;
wire n_2_10;
wire n_2_11;
wire n_2_12;
wire n_2_13;
wire n_2_14;
wire n_2_15;
wire n_2_16;
wire n_2_17;
wire n_2_18;
wire n_2_19;
wire n_2_20;
wire n_2_21;
wire n_2_22;
wire n_2_23;
wire n_2_24;
wire n_2_25;
wire n_2_26;
wire n_2_27;
wire n_2_28;
wire n_2_29;
wire n_2_30;
wire n_2_31;
wire n_2_32;
wire n_2_33;
wire n_2_34;
wire n_2_35;
wire n_2_36;
wire n_2_37;
wire n_2_38;
wire n_2_39;
wire n_2_40;
wire n_2_41;
wire n_2_42;
wire n_2_43;
wire n_2_44;
wire n_2_45;
wire n_2_46;
wire n_2_47;
wire n_2_48;
wire n_2_49;
wire n_2_50;
wire n_2_51;
wire n_2_52;
wire n_2_53;
wire n_2_54;
wire n_2_55;
wire n_2_56;
wire n_2_57;
wire n_2_58;
wire n_2_59;
wire n_2_60;
wire n_2_61;
wire n_2_62;
wire n_2_63;
wire n_2_64;
wire n_2_65;
wire n_2_66;
wire n_2_67;
wire n_2_68;
wire n_2_69;
wire n_2_70;
wire n_2_71;
wire n_2_72;
wire n_2_73;
wire n_2_74;
wire n_2_75;
wire n_2_76;
wire n_2_77;
wire n_2_78;
wire n_2_79;
wire n_2_80;
wire n_2_81;
wire n_2_82;
wire n_2_83;
wire n_2_84;
wire n_2_85;
wire n_2_86;
wire n_2_87;
wire n_2_88;
wire n_2_89;
wire n_2_90;
wire n_2_91;
wire n_2_92;
wire n_2_93;
wire n_2_94;
wire n_2_95;
wire n_2_96;
wire n_2_97;
wire n_2_98;
wire n_2_99;
wire n_2_100;
wire n_2_101;
wire n_2_102;
wire n_2_103;
wire n_2_104;
wire n_2_105;
wire n_2_106;
wire n_2_107;
wire n_2_108;
wire n_2_109;
wire n_2_110;
wire n_2_111;
wire n_2_112;
wire n_2_113;
wire n_2_114;
wire n_2_115;
wire n_2_116;
wire n_2_117;
wire n_2_118;
wire n_2_119;
wire n_2_120;
wire n_2_121;
wire n_282;
wire CTS_n_tid0_112;
wire n_281;
wire n_280;
wire n_279;
wire n_278;
wire n_277;
wire n_276;
wire n_275;
wire n_274;
wire n_273;
wire n_272;
wire n_271;
wire n_270;
wire n_269;
wire n_268;
wire n_267;
wire n_266;
wire n_265;
wire n_264;
wire n_263;
wire n_262;
wire n_261;
wire n_260;
wire n_259;
wire n_258;
wire n_257;
wire n_256;
wire n_255;
wire n_254;
wire n_253;
wire n_252;
wire n_251;
wire n_250;
wire n_249;
wire n_248;
wire n_247;
wire n_246;
wire n_245;
wire n_244;
wire n_243;
wire n_242;
wire n_241;
wire n_240;
wire n_239;
wire n_238;
wire n_237;
wire n_236;
wire n_235;
wire n_234;
wire n_233;
wire n_232;
wire n_231;
wire n_230;
wire n_229;
wire n_228;
wire n_227;
wire n_226;
wire n_225;
wire n_224;
wire n_223;
wire n_222;
wire n_221;
wire n_220;
wire n_219;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_183;
wire n_133;
wire n_216;
wire n_215;
wire n_214;
wire n_213;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_208;
wire n_207;
wire n_206;
wire n_205;
wire n_204;
wire n_203;
wire n_202;
wire n_200;
wire n_199;
wire n_198;
wire n_197;
wire n_196;
wire n_195;
wire n_194;
wire n_193;
wire n_192;
wire n_191;
wire n_190;
wire n_189;
wire n_188;
wire n_187;
wire n_186;
wire n_185;
wire n_184;
wire n_149;
wire n_182;
wire n_181;
wire n_180;
wire n_179;
wire n_178;
wire n_177;
wire n_176;
wire n_175;
wire n_174;
wire n_173;
wire n_172;
wire n_171;
wire n_170;
wire n_169;
wire n_168;
wire n_166;
wire n_165;
wire n_164;
wire n_163;
wire n_162;
wire n_161;
wire n_160;
wire n_159;
wire n_158;
wire n_157;
wire n_156;
wire n_155;
wire n_154;
wire n_153;
wire n_152;
wire n_151;
wire n_150;
wire n_218;
wire n_201;
wire n_148;
wire n_147;
wire n_146;
wire n_145;
wire n_144;
wire n_143;
wire n_66;
wire n_67;
wire n_68;
wire n_139;
wire n_138;
wire n_140;
wire n_142;
wire n_137;
wire CTS_n_tid1_16;
wire n_136;
wire n_135;
wire n_134;
wire n_132;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_127;
wire n_126;
wire n_125;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_120;
wire n_119;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_102;
wire n_141;
wire n_103;
wire n_217;
wire n_104;


INV_X1 i_2_298 (.ZN (n_2_121), .A (\count[4] ));
INV_X2 i_2_297 (.ZN (n_2_120), .A (reset));
INV_X1 i_2_296 (.ZN (n_2_119), .A (\state[2] ));
INV_X1 i_2_295 (.ZN (n_2_118), .A (\state[0] ));
XNOR2_X1 i_2_294 (.ZN (n_2_117), .A (Qbit), .B (Mbit));
NOR2_X1 i_2_293 (.ZN (n_2_116), .A1 (n_2_117), .A2 (reset));
AND2_X1 i_2_292 (.ZN (n_2_115), .A1 (n_2_120), .A2 (n_2_117));
AOI22_X1 i_2_291 (.ZN (n_2_114), .A1 (n_65), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[31] ));
INV_X1 i_2_290 (.ZN (n_282), .A (n_2_114));
AOI22_X1 i_2_289 (.ZN (n_2_113), .A1 (n_64), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[30] ));
INV_X1 i_2_288 (.ZN (n_281), .A (n_2_113));
AOI22_X1 i_2_287 (.ZN (n_2_112), .A1 (n_63), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[29] ));
INV_X1 i_2_286 (.ZN (n_280), .A (n_2_112));
AOI22_X1 i_2_285 (.ZN (n_2_111), .A1 (n_62), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[28] ));
INV_X1 i_2_284 (.ZN (n_279), .A (n_2_111));
AOI22_X1 i_2_283 (.ZN (n_2_110), .A1 (n_61), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[27] ));
INV_X1 i_2_282 (.ZN (n_278), .A (n_2_110));
AOI22_X1 i_2_281 (.ZN (n_2_109), .A1 (n_60), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[26] ));
INV_X1 i_2_280 (.ZN (n_277), .A (n_2_109));
AOI22_X1 i_2_279 (.ZN (n_2_108), .A1 (n_59), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[25] ));
INV_X1 i_2_278 (.ZN (n_276), .A (n_2_108));
AOI22_X1 i_2_277 (.ZN (n_2_107), .A1 (n_58), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[24] ));
INV_X1 i_2_276 (.ZN (n_275), .A (n_2_107));
AOI22_X1 i_2_275 (.ZN (n_2_106), .A1 (n_57), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[23] ));
INV_X1 i_2_274 (.ZN (n_274), .A (n_2_106));
AOI22_X1 i_2_273 (.ZN (n_2_105), .A1 (n_56), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[22] ));
INV_X1 i_2_272 (.ZN (n_273), .A (n_2_105));
AOI22_X1 i_2_271 (.ZN (n_2_104), .A1 (n_55), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[21] ));
INV_X1 i_2_270 (.ZN (n_272), .A (n_2_104));
AOI22_X1 i_2_269 (.ZN (n_2_103), .A1 (n_54), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[20] ));
INV_X1 i_2_268 (.ZN (n_271), .A (n_2_103));
AOI22_X1 i_2_267 (.ZN (n_2_102), .A1 (n_53), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[19] ));
INV_X1 i_2_266 (.ZN (n_270), .A (n_2_102));
AOI22_X1 i_2_265 (.ZN (n_2_101), .A1 (n_52), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[18] ));
INV_X1 i_2_264 (.ZN (n_269), .A (n_2_101));
AOI22_X1 i_2_263 (.ZN (n_2_100), .A1 (n_51), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[17] ));
INV_X1 i_2_262 (.ZN (n_268), .A (n_2_100));
AOI22_X1 i_2_261 (.ZN (n_2_99), .A1 (n_50), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[16] ));
INV_X1 i_2_260 (.ZN (n_267), .A (n_2_99));
AOI22_X1 i_2_259 (.ZN (n_2_98), .A1 (n_49), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[15] ));
INV_X1 i_2_258 (.ZN (n_266), .A (n_2_98));
AOI22_X1 i_2_257 (.ZN (n_2_97), .A1 (n_48), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[14] ));
INV_X1 i_2_256 (.ZN (n_265), .A (n_2_97));
AOI22_X1 i_2_255 (.ZN (n_2_96), .A1 (n_47), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[13] ));
INV_X1 i_2_254 (.ZN (n_264), .A (n_2_96));
AOI22_X1 i_2_253 (.ZN (n_2_95), .A1 (n_46), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[12] ));
INV_X1 i_2_252 (.ZN (n_263), .A (n_2_95));
AOI22_X1 i_2_251 (.ZN (n_2_94), .A1 (n_45), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[11] ));
INV_X1 i_2_250 (.ZN (n_262), .A (n_2_94));
AOI22_X1 i_2_249 (.ZN (n_2_93), .A1 (n_44), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[10] ));
INV_X1 i_2_248 (.ZN (n_261), .A (n_2_93));
AOI22_X1 i_2_247 (.ZN (n_2_92), .A1 (n_43), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[9] ));
INV_X1 i_2_246 (.ZN (n_260), .A (n_2_92));
AOI22_X1 i_2_245 (.ZN (n_2_91), .A1 (n_42), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[8] ));
INV_X1 i_2_244 (.ZN (n_259), .A (n_2_91));
AOI22_X1 i_2_243 (.ZN (n_2_90), .A1 (n_41), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[7] ));
INV_X1 i_2_242 (.ZN (n_258), .A (n_2_90));
AOI22_X1 i_2_241 (.ZN (n_2_89), .A1 (n_40), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[6] ));
INV_X1 i_2_240 (.ZN (n_257), .A (n_2_89));
AOI22_X1 i_2_239 (.ZN (n_2_88), .A1 (n_39), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[5] ));
INV_X1 i_2_238 (.ZN (n_256), .A (n_2_88));
AOI22_X1 i_2_237 (.ZN (n_2_87), .A1 (n_38), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[4] ));
INV_X1 i_2_236 (.ZN (n_255), .A (n_2_87));
AOI22_X1 i_2_235 (.ZN (n_2_86), .A1 (n_37), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[3] ));
INV_X1 i_2_234 (.ZN (n_254), .A (n_2_86));
AOI22_X1 i_2_233 (.ZN (n_2_85), .A1 (n_36), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[2] ));
INV_X1 i_2_232 (.ZN (n_253), .A (n_2_85));
AOI22_X1 i_2_231 (.ZN (n_2_84), .A1 (n_35), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\Acc[1] ));
INV_X1 i_2_230 (.ZN (n_252), .A (n_2_84));
AOI22_X1 i_2_229 (.ZN (n_2_83), .A1 (n_34), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\Acc[0] ));
INV_X1 i_2_228 (.ZN (n_251), .A (n_2_83));
AOI22_X1 i_2_227 (.ZN (n_2_82), .A1 (n_33), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[31] ));
INV_X1 i_2_226 (.ZN (n_250), .A (n_2_82));
AOI22_X1 i_2_225 (.ZN (n_2_81), .A1 (n_32), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[30] ));
INV_X1 i_2_224 (.ZN (n_249), .A (n_2_81));
AOI22_X1 i_2_223 (.ZN (n_2_80), .A1 (n_31), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[29] ));
INV_X1 i_2_222 (.ZN (n_248), .A (n_2_80));
AOI22_X1 i_2_221 (.ZN (n_2_79), .A1 (n_30), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[28] ));
INV_X1 i_2_220 (.ZN (n_247), .A (n_2_79));
AOI22_X1 i_2_219 (.ZN (n_2_78), .A1 (n_29), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[27] ));
INV_X1 i_2_218 (.ZN (n_246), .A (n_2_78));
AOI22_X1 i_2_217 (.ZN (n_2_77), .A1 (n_28), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[26] ));
INV_X1 i_2_216 (.ZN (n_245), .A (n_2_77));
AOI22_X1 i_2_215 (.ZN (n_2_76), .A1 (n_27), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[25] ));
INV_X1 i_2_214 (.ZN (n_244), .A (n_2_76));
AOI22_X1 i_2_213 (.ZN (n_2_75), .A1 (n_26), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[24] ));
INV_X1 i_2_212 (.ZN (n_243), .A (n_2_75));
AOI22_X1 i_2_211 (.ZN (n_2_74), .A1 (n_25), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[23] ));
INV_X1 i_2_210 (.ZN (n_242), .A (n_2_74));
AOI22_X1 i_2_209 (.ZN (n_2_73), .A1 (n_24), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[22] ));
INV_X1 i_2_208 (.ZN (n_241), .A (n_2_73));
AOI22_X1 i_2_207 (.ZN (n_2_72), .A1 (n_23), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[21] ));
INV_X1 i_2_206 (.ZN (n_240), .A (n_2_72));
AOI22_X1 i_2_205 (.ZN (n_2_71), .A1 (n_22), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[20] ));
INV_X1 i_2_204 (.ZN (n_239), .A (n_2_71));
AOI22_X1 i_2_203 (.ZN (n_2_70), .A1 (n_21), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[19] ));
INV_X1 i_2_202 (.ZN (n_238), .A (n_2_70));
AOI22_X1 i_2_201 (.ZN (n_2_69), .A1 (n_20), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[18] ));
INV_X1 i_2_200 (.ZN (n_237), .A (n_2_69));
AOI22_X1 i_2_199 (.ZN (n_2_68), .A1 (n_19), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[17] ));
INV_X1 i_2_198 (.ZN (n_236), .A (n_2_68));
AOI22_X1 i_2_197 (.ZN (n_2_67), .A1 (n_18), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[16] ));
INV_X1 i_2_196 (.ZN (n_235), .A (n_2_67));
AOI22_X1 i_2_195 (.ZN (n_2_66), .A1 (n_17), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[15] ));
INV_X1 i_2_194 (.ZN (n_234), .A (n_2_66));
AOI22_X1 i_2_193 (.ZN (n_2_65), .A1 (n_16), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[14] ));
INV_X1 i_2_192 (.ZN (n_233), .A (n_2_65));
AOI22_X1 i_2_191 (.ZN (n_2_64), .A1 (n_15), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[13] ));
INV_X1 i_2_190 (.ZN (n_232), .A (n_2_64));
AOI22_X1 i_2_189 (.ZN (n_2_63), .A1 (n_14), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[12] ));
INV_X1 i_2_188 (.ZN (n_231), .A (n_2_63));
AOI22_X1 i_2_187 (.ZN (n_2_62), .A1 (n_13), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[11] ));
INV_X1 i_2_186 (.ZN (n_230), .A (n_2_62));
AOI22_X1 i_2_185 (.ZN (n_2_61), .A1 (n_12), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[10] ));
INV_X1 i_2_184 (.ZN (n_229), .A (n_2_61));
AOI22_X1 i_2_183 (.ZN (n_2_60), .A1 (n_11), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[9] ));
INV_X1 i_2_182 (.ZN (n_228), .A (n_2_60));
AOI22_X1 i_2_181 (.ZN (n_2_59), .A1 (n_10), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[8] ));
INV_X1 i_2_180 (.ZN (n_227), .A (n_2_59));
AOI22_X1 i_2_179 (.ZN (n_2_58), .A1 (n_9), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[7] ));
INV_X1 i_2_178 (.ZN (n_226), .A (n_2_58));
AOI22_X1 i_2_177 (.ZN (n_2_57), .A1 (n_8), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[6] ));
INV_X1 i_2_176 (.ZN (n_225), .A (n_2_57));
AOI22_X1 i_2_175 (.ZN (n_2_56), .A1 (n_7), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[5] ));
INV_X1 i_2_174 (.ZN (n_224), .A (n_2_56));
AOI22_X1 i_2_173 (.ZN (n_2_55), .A1 (n_6), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[4] ));
INV_X1 i_2_172 (.ZN (n_223), .A (n_2_55));
AOI22_X1 i_2_171 (.ZN (n_2_54), .A1 (n_5), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[3] ));
INV_X1 i_2_170 (.ZN (n_222), .A (n_2_54));
AOI22_X1 i_2_169 (.ZN (n_2_53), .A1 (n_4), .A2 (hfn_ipo_n11), .B1 (hfn_ipo_n9), .B2 (\inputQ_reg[2] ));
INV_X1 i_2_168 (.ZN (n_221), .A (n_2_53));
AOI22_X1 i_2_167 (.ZN (n_2_52), .A1 (n_3), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[1] ));
INV_X1 i_2_166 (.ZN (n_220), .A (n_2_52));
AOI22_X1 i_2_165 (.ZN (n_2_51), .A1 (n_2), .A2 (hfn_ipo_n12), .B1 (hfn_ipo_n10), .B2 (\inputQ_reg[0] ));
INV_X1 i_2_164 (.ZN (n_219), .A (n_2_51));
OR3_X1 i_2_163 (.ZN (n_2_50), .A1 (n_2_118), .A2 (\state[1] ), .A3 (\state[2] ));
NAND2_X1 i_2_162 (.ZN (n_218), .A1 (n_2_120), .A2 (n_2_50));
NOR2_X1 i_2_161 (.ZN (n_2_49), .A1 (\count[5] ), .A2 (reset));
OR2_X1 i_2_160 (.ZN (n_2_48), .A1 (\count[5] ), .A2 (reset));
AOI21_X1 i_2_159 (.ZN (n_217), .A (n_2_49), .B1 (n_2_50), .B2 (n_2_120));
NOR2_X1 i_2_158 (.ZN (n_2_47), .A1 (\state[1] ), .A2 (\state[0] ));
INV_X1 i_2_157 (.ZN (n_2_46), .A (n_2_47));
NAND2_X2 i_2_156 (.ZN (n_2_45), .A1 (n_2_47), .A2 (n_2_119));
MUX2_X1 i_2_155 (.Z (n_2_44), .A (\Acc[0] ), .B (\add_output[0] ), .S (lsb_reg));
MUX2_X1 i_2_154 (.Z (n_216), .A (inputQ_wire[31]), .B (n_2_44), .S (n_2_45));
MUX2_X1 i_2_153 (.Z (n_215), .A (inputQ_wire[30]), .B (\inputQ_reg[31] ), .S (n_2_45));
MUX2_X1 i_2_152 (.Z (n_214), .A (inputQ_wire[29]), .B (\inputQ_reg[30] ), .S (n_2_45));
MUX2_X1 i_2_151 (.Z (n_213), .A (inputQ_wire[28]), .B (\inputQ_reg[29] ), .S (n_2_45));
MUX2_X1 i_2_150 (.Z (n_212), .A (inputQ_wire[27]), .B (\inputQ_reg[28] ), .S (n_2_45));
MUX2_X1 i_2_149 (.Z (n_211), .A (inputQ_wire[26]), .B (\inputQ_reg[27] ), .S (n_2_45));
MUX2_X1 i_2_148 (.Z (n_210), .A (inputQ_wire[25]), .B (\inputQ_reg[26] ), .S (n_2_45));
MUX2_X1 i_2_147 (.Z (n_209), .A (inputQ_wire[24]), .B (\inputQ_reg[25] ), .S (n_2_45));
MUX2_X1 i_2_146 (.Z (n_208), .A (inputQ_wire[23]), .B (\inputQ_reg[24] ), .S (n_2_45));
MUX2_X1 i_2_145 (.Z (n_207), .A (inputQ_wire[22]), .B (\inputQ_reg[23] ), .S (n_2_45));
MUX2_X1 i_2_144 (.Z (n_206), .A (inputQ_wire[21]), .B (\inputQ_reg[22] ), .S (n_2_45));
MUX2_X1 i_2_143 (.Z (n_205), .A (inputQ_wire[20]), .B (\inputQ_reg[21] ), .S (n_2_45));
MUX2_X1 i_2_142 (.Z (n_204), .A (inputQ_wire[19]), .B (\inputQ_reg[20] ), .S (n_2_45));
MUX2_X1 i_2_141 (.Z (n_203), .A (inputQ_wire[18]), .B (\inputQ_reg[19] ), .S (n_2_45));
MUX2_X1 i_2_140 (.Z (n_202), .A (inputQ_wire[17]), .B (\inputQ_reg[18] ), .S (n_2_45));
MUX2_X1 i_2_139 (.Z (n_200), .A (inputQ_wire[16]), .B (\inputQ_reg[17] ), .S (n_2_45));
MUX2_X1 i_2_138 (.Z (n_199), .A (inputQ_wire[15]), .B (\inputQ_reg[16] ), .S (n_2_45));
MUX2_X1 i_2_137 (.Z (n_198), .A (inputQ_wire[14]), .B (\inputQ_reg[15] ), .S (n_2_45));
MUX2_X1 i_2_136 (.Z (n_197), .A (inputQ_wire[13]), .B (\inputQ_reg[14] ), .S (n_2_45));
MUX2_X1 i_2_135 (.Z (n_196), .A (inputQ_wire[12]), .B (\inputQ_reg[13] ), .S (n_2_45));
MUX2_X1 i_2_134 (.Z (n_195), .A (inputQ_wire[11]), .B (\inputQ_reg[12] ), .S (n_2_45));
MUX2_X1 i_2_133 (.Z (n_194), .A (inputQ_wire[10]), .B (\inputQ_reg[11] ), .S (n_2_45));
MUX2_X1 i_2_132 (.Z (n_193), .A (inputQ_wire[9]), .B (\inputQ_reg[10] ), .S (n_2_45));
MUX2_X1 i_2_131 (.Z (n_192), .A (inputQ_wire[8]), .B (\inputQ_reg[9] ), .S (n_2_45));
MUX2_X1 i_2_130 (.Z (n_191), .A (inputQ_wire[7]), .B (\inputQ_reg[8] ), .S (n_2_45));
MUX2_X1 i_2_129 (.Z (n_190), .A (inputQ_wire[6]), .B (\inputQ_reg[7] ), .S (n_2_45));
MUX2_X1 i_2_128 (.Z (n_189), .A (inputQ_wire[5]), .B (\inputQ_reg[6] ), .S (n_2_45));
MUX2_X1 i_2_127 (.Z (n_188), .A (inputQ_wire[4]), .B (\inputQ_reg[5] ), .S (n_2_45));
MUX2_X1 i_2_126 (.Z (n_187), .A (inputQ_wire[3]), .B (\inputQ_reg[4] ), .S (n_2_45));
MUX2_X1 i_2_125 (.Z (n_186), .A (inputQ_wire[2]), .B (\inputQ_reg[3] ), .S (n_2_45));
MUX2_X1 i_2_124 (.Z (n_185), .A (inputQ_wire[1]), .B (\inputQ_reg[2] ), .S (n_2_45));
MUX2_X1 i_2_123 (.Z (n_184), .A (inputQ_wire[0]), .B (\inputQ_reg[1] ), .S (n_2_45));
NOR2_X1 i_2_122 (.ZN (n_183), .A1 (n_2_46), .A2 (reset));
AND2_X2 i_2_121 (.ZN (n_2_43), .A1 (n_2_120), .A2 (lsb_reg));
NAND2_X1 i_2_120 (.ZN (n_2_42), .A1 (n_2_120), .A2 (lsb_reg));
AND2_X1 i_2_119 (.ZN (n_182), .A1 (c_output), .A2 (n_2_43));
NOR2_X4 i_2_118 (.ZN (n_2_41), .A1 (reset), .A2 (lsb_reg));
AOI22_X1 i_2_117 (.ZN (n_2_40), .A1 (\add_output[31] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[31] ));
INV_X1 i_2_116 (.ZN (n_181), .A (n_2_40));
AOI22_X1 i_2_115 (.ZN (n_2_39), .A1 (\add_output[30] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[30] ));
INV_X1 i_2_114 (.ZN (n_180), .A (n_2_39));
AOI22_X1 i_2_113 (.ZN (n_2_38), .A1 (\add_output[29] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[29] ));
INV_X1 i_2_112 (.ZN (n_179), .A (n_2_38));
AOI22_X1 i_2_111 (.ZN (n_2_37), .A1 (\add_output[28] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[28] ));
INV_X1 i_2_110 (.ZN (n_178), .A (n_2_37));
AOI22_X1 i_2_109 (.ZN (n_2_36), .A1 (\add_output[27] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[27] ));
INV_X1 i_2_108 (.ZN (n_177), .A (n_2_36));
AOI22_X1 i_2_107 (.ZN (n_2_35), .A1 (\add_output[26] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[26] ));
INV_X1 i_2_106 (.ZN (n_176), .A (n_2_35));
AOI22_X1 i_2_105 (.ZN (n_2_34), .A1 (\add_output[25] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[25] ));
INV_X1 i_2_104 (.ZN (n_175), .A (n_2_34));
AOI22_X1 i_2_103 (.ZN (n_2_33), .A1 (\add_output[24] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[24] ));
INV_X1 i_2_102 (.ZN (n_174), .A (n_2_33));
AOI22_X1 i_2_101 (.ZN (n_2_32), .A1 (\add_output[23] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[23] ));
INV_X1 i_2_100 (.ZN (n_173), .A (n_2_32));
AOI22_X1 i_2_99 (.ZN (n_2_31), .A1 (\add_output[22] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[22] ));
INV_X1 i_2_98 (.ZN (n_172), .A (n_2_31));
AOI22_X1 i_2_97 (.ZN (n_2_30), .A1 (\add_output[21] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[21] ));
INV_X1 i_2_96 (.ZN (n_171), .A (n_2_30));
AOI22_X1 i_2_95 (.ZN (n_2_29), .A1 (\add_output[20] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[20] ));
INV_X1 i_2_94 (.ZN (n_170), .A (n_2_29));
AOI22_X1 i_2_93 (.ZN (n_2_28), .A1 (\add_output[19] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[19] ));
INV_X1 i_2_92 (.ZN (n_169), .A (n_2_28));
AOI22_X1 i_2_91 (.ZN (n_2_27), .A1 (\add_output[18] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[18] ));
INV_X1 i_2_90 (.ZN (n_168), .A (n_2_27));
AOI22_X1 i_2_89 (.ZN (n_2_26), .A1 (\add_output[17] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[17] ));
INV_X1 i_2_88 (.ZN (n_166), .A (n_2_26));
AOI22_X1 i_2_87 (.ZN (n_2_25), .A1 (\add_output[16] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[16] ));
INV_X1 i_2_86 (.ZN (n_165), .A (n_2_25));
AOI22_X1 i_2_85 (.ZN (n_2_24), .A1 (\add_output[15] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[15] ));
INV_X1 i_2_84 (.ZN (n_164), .A (n_2_24));
AOI22_X1 i_2_83 (.ZN (n_2_23), .A1 (\add_output[14] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[14] ));
INV_X1 i_2_82 (.ZN (n_163), .A (n_2_23));
AOI22_X1 i_2_81 (.ZN (n_2_22), .A1 (\add_output[13] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[13] ));
INV_X1 i_2_80 (.ZN (n_162), .A (n_2_22));
AOI22_X1 i_2_79 (.ZN (n_2_21), .A1 (\add_output[12] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[12] ));
INV_X1 i_2_78 (.ZN (n_161), .A (n_2_21));
AOI22_X1 i_2_77 (.ZN (n_2_20), .A1 (\add_output[11] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[11] ));
INV_X1 i_2_76 (.ZN (n_160), .A (n_2_20));
AOI22_X1 i_2_75 (.ZN (n_2_19), .A1 (\add_output[10] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[10] ));
INV_X1 i_2_74 (.ZN (n_159), .A (n_2_19));
AOI22_X1 i_2_73 (.ZN (n_2_18), .A1 (\add_output[9] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[9] ));
INV_X1 i_2_72 (.ZN (n_158), .A (n_2_18));
AOI22_X1 i_2_71 (.ZN (n_2_17), .A1 (\add_output[8] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[8] ));
INV_X1 i_2_70 (.ZN (n_157), .A (n_2_17));
AOI22_X1 i_2_69 (.ZN (n_2_16), .A1 (\add_output[7] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[7] ));
INV_X1 i_2_68 (.ZN (n_156), .A (n_2_16));
AOI22_X1 i_2_67 (.ZN (n_2_15), .A1 (\add_output[6] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[6] ));
INV_X1 i_2_66 (.ZN (n_155), .A (n_2_15));
AOI22_X1 i_2_65 (.ZN (n_2_14), .A1 (\add_output[5] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[5] ));
INV_X1 i_2_64 (.ZN (n_154), .A (n_2_14));
AOI22_X1 i_2_63 (.ZN (n_2_13), .A1 (\add_output[4] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[4] ));
INV_X1 i_2_62 (.ZN (n_153), .A (n_2_13));
AOI22_X1 i_2_61 (.ZN (n_2_12), .A1 (\add_output[3] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[3] ));
INV_X1 i_2_60 (.ZN (n_152), .A (n_2_12));
AOI22_X1 i_2_59 (.ZN (n_2_11), .A1 (\add_output[2] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[2] ));
INV_X1 i_2_58 (.ZN (n_151), .A (n_2_11));
AOI22_X1 i_2_57 (.ZN (n_2_10), .A1 (\add_output[1] ), .A2 (n_2_43), .B1 (n_2_41), .B2 (\Acc[1] ));
INV_X1 i_2_56 (.ZN (n_150), .A (n_2_10));
AOI21_X1 i_2_55 (.ZN (n_2_9), .A (reset), .B1 (\state[2] ), .B2 (n_2_47));
INV_X1 i_2_54 (.ZN (n_149), .A (n_2_9));
AND3_X1 i_2_53 (.ZN (n_2_8), .A1 (\count[2] ), .A2 (\count[1] ), .A3 (\count[0] ));
NAND2_X1 i_2_52 (.ZN (n_2_7), .A1 (\count[3] ), .A2 (n_2_8));
NOR3_X1 i_2_51 (.ZN (n_148), .A1 (n_2_121), .A2 (n_2_48), .A3 (n_2_7));
NAND2_X1 i_2_50 (.ZN (n_2_6), .A1 (n_2_49), .A2 (n_2_121));
NAND3_X1 i_2_49 (.ZN (n_2_5), .A1 (n_2_7), .A2 (n_2_49), .A3 (\count[4] ));
OAI21_X1 i_2_48 (.ZN (n_147), .A (n_2_5), .B1 (n_2_6), .B2 (n_2_7));
OAI21_X1 i_2_47 (.ZN (n_2_4), .A (n_2_49), .B1 (n_2_8), .B2 (\count[3] ));
AOI21_X1 i_2_46 (.ZN (n_146), .A (n_2_4), .B1 (n_2_8), .B2 (\count[3] ));
AOI21_X1 i_2_45 (.ZN (n_2_3), .A (\count[2] ), .B1 (\count[1] ), .B2 (\count[0] ));
NOR3_X1 i_2_44 (.ZN (n_145), .A1 (n_2_48), .A2 (n_2_8), .A3 (n_2_3));
OAI21_X1 i_2_43 (.ZN (n_2_2), .A (n_2_49), .B1 (\count[0] ), .B2 (\count[1] ));
AOI21_X1 i_2_42 (.ZN (n_144), .A (n_2_2), .B1 (\count[0] ), .B2 (\count[1] ));
NOR2_X1 i_2_41 (.ZN (n_143), .A1 (n_2_48), .A2 (\count[0] ));
NAND2_X1 i_2_40 (.ZN (n_2_1), .A1 (n_2_119), .A2 (\state[1] ));
AOI211_X1 i_2_39 (.ZN (n_142), .A (reset), .B (n_2_1), .C1 (lsb_reg), .C2 (n_2_118));
NOR2_X1 i_2_38 (.ZN (n_141), .A1 (n_2_50), .A2 (n_2_48));
OAI33_X1 i_2_37 (.ZN (n_140), .A1 (n_2_50), .A2 (reset), .A3 (\count[5] ), .B1 (\state[0] )
    , .B2 (n_2_42), .B3 (n_2_1));
NOR2_X1 i_2_36 (.ZN (n_2_0), .A1 (\state[2] ), .A2 (start));
OAI33_X1 i_2_35 (.ZN (n_139), .A1 (reset), .A2 (n_2_46), .A3 (n_2_0), .B1 (n_2_1)
    , .B2 (n_2_42), .B3 (\state[0] ));
NAND3_X1 i_2_34 (.ZN (n_138), .A1 (n_2_120), .A2 (n_2_46), .A3 (\state[2] ));
AND2_X1 i_2_33 (.ZN (n_137), .A1 (n_2_120), .A2 (n_100));
AND2_X1 i_2_32 (.ZN (n_136), .A1 (n_2_120), .A2 (n_99));
AND2_X1 i_2_31 (.ZN (n_135), .A1 (n_2_120), .A2 (n_98));
AND2_X1 i_2_30 (.ZN (n_134), .A1 (n_2_120), .A2 (n_97));
AND2_X1 i_2_29 (.ZN (n_132), .A1 (n_2_120), .A2 (n_96));
AND2_X1 i_2_28 (.ZN (n_131), .A1 (n_2_120), .A2 (n_95));
AND2_X1 i_2_27 (.ZN (n_130), .A1 (n_2_120), .A2 (n_94));
AND2_X1 i_2_26 (.ZN (n_129), .A1 (n_2_120), .A2 (n_93));
AND2_X1 i_2_25 (.ZN (n_128), .A1 (n_2_120), .A2 (n_92));
AND2_X1 i_2_24 (.ZN (n_127), .A1 (n_2_120), .A2 (n_91));
AND2_X1 i_2_23 (.ZN (n_126), .A1 (n_2_120), .A2 (n_90));
AND2_X1 i_2_22 (.ZN (n_125), .A1 (n_2_120), .A2 (n_89));
AND2_X1 i_2_21 (.ZN (n_124), .A1 (n_2_120), .A2 (n_88));
AND2_X1 i_2_20 (.ZN (n_123), .A1 (n_2_120), .A2 (n_87));
AND2_X1 i_2_19 (.ZN (n_122), .A1 (n_2_120), .A2 (n_86));
AND2_X1 i_2_18 (.ZN (n_121), .A1 (n_2_120), .A2 (n_85));
AND2_X1 i_2_17 (.ZN (n_120), .A1 (n_2_120), .A2 (n_84));
AND2_X1 i_2_16 (.ZN (n_119), .A1 (n_2_120), .A2 (n_83));
AND2_X1 i_2_15 (.ZN (n_118), .A1 (n_2_120), .A2 (n_82));
AND2_X1 i_2_14 (.ZN (n_117), .A1 (n_2_120), .A2 (n_81));
AND2_X1 i_2_13 (.ZN (n_116), .A1 (n_2_120), .A2 (n_80));
AND2_X1 i_2_12 (.ZN (n_115), .A1 (n_2_120), .A2 (n_79));
AND2_X1 i_2_11 (.ZN (n_114), .A1 (n_2_120), .A2 (n_78));
AND2_X1 i_2_10 (.ZN (n_113), .A1 (n_2_120), .A2 (n_77));
AND2_X1 i_2_9 (.ZN (n_112), .A1 (n_2_120), .A2 (n_76));
AND2_X1 i_2_8 (.ZN (n_111), .A1 (n_2_120), .A2 (n_75));
AND2_X1 i_2_7 (.ZN (n_110), .A1 (n_2_120), .A2 (n_74));
AND2_X1 i_2_6 (.ZN (n_109), .A1 (n_2_120), .A2 (n_73));
AND2_X1 i_2_5 (.ZN (n_108), .A1 (n_2_120), .A2 (n_72));
AND2_X1 i_2_4 (.ZN (n_107), .A1 (n_2_120), .A2 (n_71));
AND2_X1 i_2_3 (.ZN (n_106), .A1 (n_2_120), .A2 (n_70));
AND2_X1 i_2_2 (.ZN (n_105), .A1 (n_2_120), .A2 (n_69));
OAI21_X1 i_2_1 (.ZN (n_104), .A (n_2_120), .B1 (n_2_118), .B2 (n_2_1));
AND2_X1 i_2_0 (.ZN (n_103), .A1 (n_2_120), .A2 (n_101));
CLKGATETST_X8 clk_gate_c_output_reg (.GCK (CTS_n_tid1_17), .CK (CTS_n_tid0_209), .E (n_104), .SE (1'b0 ));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid0_188), .CK (CTS_n_tid0_209), .E (n_217), .SE (1'b0 ));
DFF_X1 start_reg (.Q (start), .CK (CTS_n_tid0_121), .D (reset));
DFF_X1 c_output_reg (.Q (c_output), .CK (CTS_n_tid1_16), .D (n_103));
MUX2_X1 lsb_reg_reg_enable_mux_0 (.Z (n_102), .A (lsb_reg), .B (\inputQ_reg[0] ), .S (n_141));
DFF_X1 lsb_reg_reg (.Q (lsb_reg), .CK (CTS_n_tid0_198), .D (n_102));
datapath__0_17 i_16 (.p_0 ({n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, 
    n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, 
    n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69}), .Acc ({\Acc[31] , 
    \Acc[30] , \Acc[29] , \Acc[28] , \Acc[27] , \Acc[26] , \Acc[25] , \Acc[24] , 
    \Acc[23] , \Acc[22] , \Acc[21] , \Acc[20] , \Acc[19] , \Acc[18] , \Acc[17] , 
    \Acc[16] , \Acc[15] , \Acc[14] , \Acc[13] , \Acc[12] , \Acc[11] , \Acc[10] , 
    \Acc[9] , \Acc[8] , \Acc[7] , \Acc[6] , \Acc[5] , \Acc[4] , \Acc[3] , \Acc[2] , 
    \Acc[1] , \Acc[0] }), .inputM_wire ({inputM_wire[31], inputM_wire[30], inputM_wire[29], 
    inputM_wire[28], inputM_wire[27], inputM_wire[26], inputM_wire[25], inputM_wire[24], 
    inputM_wire[23], inputM_wire[22], inputM_wire[21], inputM_wire[20], inputM_wire[19], 
    inputM_wire[18], inputM_wire[17], inputM_wire[16], inputM_wire[15], inputM_wire[14], 
    inputM_wire[13], inputM_wire[12], inputM_wire[11], inputM_wire[10], inputM_wire[9], 
    inputM_wire[8], inputM_wire[7], inputM_wire[6], inputM_wire[5], inputM_wire[4], 
    inputM_wire[3], inputM_wire[2], inputM_wire[1], inputM_wire[0]}));
DFF_X1 \add_output_reg[0]  (.Q (\add_output[0] ), .CK (CTS_n_tid1_16), .D (n_105));
DFF_X1 \add_output_reg[1]  (.Q (\add_output[1] ), .CK (CTS_n_tid1_16), .D (n_106));
DFF_X1 \add_output_reg[2]  (.Q (\add_output[2] ), .CK (CTS_n_tid1_16), .D (n_107));
DFF_X1 \add_output_reg[3]  (.Q (\add_output[3] ), .CK (CTS_n_tid1_16), .D (n_108));
DFF_X1 \add_output_reg[4]  (.Q (\add_output[4] ), .CK (CTS_n_tid1_16), .D (n_109));
DFF_X1 \add_output_reg[5]  (.Q (\add_output[5] ), .CK (CTS_n_tid1_16), .D (n_110));
DFF_X1 \add_output_reg[6]  (.Q (\add_output[6] ), .CK (CTS_n_tid1_16), .D (n_111));
DFF_X1 \add_output_reg[7]  (.Q (\add_output[7] ), .CK (CTS_n_tid1_16), .D (n_112));
DFF_X1 \add_output_reg[8]  (.Q (\add_output[8] ), .CK (CTS_n_tid1_16), .D (n_113));
DFF_X1 \add_output_reg[9]  (.Q (\add_output[9] ), .CK (CTS_n_tid1_16), .D (n_114));
DFF_X1 \add_output_reg[10]  (.Q (\add_output[10] ), .CK (CTS_n_tid1_16), .D (n_115));
DFF_X1 \add_output_reg[11]  (.Q (\add_output[11] ), .CK (CTS_n_tid1_16), .D (n_116));
DFF_X1 \add_output_reg[12]  (.Q (\add_output[12] ), .CK (CTS_n_tid1_16), .D (n_117));
DFF_X1 \add_output_reg[13]  (.Q (\add_output[13] ), .CK (CTS_n_tid1_16), .D (n_118));
DFF_X1 \add_output_reg[14]  (.Q (\add_output[14] ), .CK (CTS_n_tid1_16), .D (n_119));
DFF_X1 \add_output_reg[15]  (.Q (\add_output[15] ), .CK (CTS_n_tid1_16), .D (n_120));
DFF_X1 \add_output_reg[16]  (.Q (\add_output[16] ), .CK (CTS_n_tid1_16), .D (n_121));
DFF_X1 \add_output_reg[17]  (.Q (\add_output[17] ), .CK (CTS_n_tid1_16), .D (n_122));
DFF_X1 \add_output_reg[18]  (.Q (\add_output[18] ), .CK (CTS_n_tid1_16), .D (n_123));
DFF_X1 \add_output_reg[19]  (.Q (\add_output[19] ), .CK (CTS_n_tid1_16), .D (n_124));
DFF_X1 \add_output_reg[20]  (.Q (\add_output[20] ), .CK (CTS_n_tid1_16), .D (n_125));
DFF_X1 \add_output_reg[21]  (.Q (\add_output[21] ), .CK (CTS_n_tid1_16), .D (n_126));
DFF_X1 \add_output_reg[22]  (.Q (\add_output[22] ), .CK (CTS_n_tid1_16), .D (n_127));
DFF_X1 \add_output_reg[23]  (.Q (\add_output[23] ), .CK (CTS_n_tid1_16), .D (n_128));
DFF_X1 \add_output_reg[24]  (.Q (\add_output[24] ), .CK (CTS_n_tid1_16), .D (n_129));
DFF_X1 \add_output_reg[25]  (.Q (\add_output[25] ), .CK (CTS_n_tid1_16), .D (n_130));
DFF_X1 \add_output_reg[26]  (.Q (\add_output[26] ), .CK (CTS_n_tid1_16), .D (n_131));
DFF_X1 \add_output_reg[27]  (.Q (\add_output[27] ), .CK (CTS_n_tid1_16), .D (n_132));
DFF_X1 \add_output_reg[28]  (.Q (\add_output[28] ), .CK (CTS_n_tid1_16), .D (n_134));
DFF_X1 \add_output_reg[29]  (.Q (\add_output[29] ), .CK (CTS_n_tid1_16), .D (n_135));
DFF_X1 \add_output_reg[30]  (.Q (\add_output[30] ), .CK (CTS_n_tid1_16), .D (n_136));
DFF_X1 \add_output_reg[31]  (.Q (\add_output[31] ), .CK (CTS_n_tid1_16), .D (n_137));
MUX2_X1 i_1_2 (.Z (n_68), .A (\state[2] ), .B (n_142), .S (n_138));
MUX2_X1 i_1_1 (.Z (n_67), .A (\state[1] ), .B (n_140), .S (n_138));
MUX2_X1 i_1_0 (.Z (n_66), .A (\state[0] ), .B (n_139), .S (n_138));
DFF_X1 \state_reg[2]  (.Q (\state[2] ), .CK (CTS_n_tid0_198), .D (n_68));
DFF_X1 \state_reg[1]  (.Q (\state[1] ), .CK (CTS_n_tid0_198), .D (n_67));
DFF_X1 \state_reg[0]  (.Q (\state[0] ), .CK (CTS_n_tid0_198), .D (n_66));
DFF_X1 \count_reg[0]  (.Q (\count[0] ), .CK (n_201), .D (n_143));
DFF_X1 \count_reg[1]  (.Q (\count[1] ), .CK (n_201), .D (n_144));
DFF_X1 \count_reg[2]  (.Q (\count[2] ), .CK (n_201), .D (n_145));
DFF_X1 \count_reg[3]  (.Q (\count[3] ), .CK (n_201), .D (n_146));
DFF_X1 \count_reg[4]  (.Q (\count[4] ), .CK (n_201), .D (n_147));
DFF_X1 \count_reg[5]  (.Q (\count[5] ), .CK (n_201), .D (n_148));
CLKGATETST_X1 clk_gate_count_reg (.GCK (n_201), .CK (CTS_n_tid0_209), .E (n_218), .SE (1'b0 ));
DFF_X1 \Acc_reg[0]  (.Q (\Acc[0] ), .CK (CTS_n_tid0_49), .D (n_150));
DFF_X1 \Acc_reg[1]  (.Q (\Acc[1] ), .CK (CTS_n_tid0_49), .D (n_151));
DFF_X1 \Acc_reg[2]  (.Q (\Acc[2] ), .CK (CTS_n_tid0_49), .D (n_152));
DFF_X1 \Acc_reg[3]  (.Q (\Acc[3] ), .CK (CTS_n_tid0_49), .D (n_153));
DFF_X1 \Acc_reg[4]  (.Q (\Acc[4] ), .CK (CTS_n_tid0_49), .D (n_154));
DFF_X1 \Acc_reg[5]  (.Q (\Acc[5] ), .CK (CTS_n_tid0_49), .D (n_155));
DFF_X1 \Acc_reg[6]  (.Q (\Acc[6] ), .CK (CTS_n_tid0_49), .D (n_156));
DFF_X1 \Acc_reg[7]  (.Q (\Acc[7] ), .CK (CTS_n_tid0_49), .D (n_157));
DFF_X1 \Acc_reg[8]  (.Q (\Acc[8] ), .CK (CTS_n_tid0_49), .D (n_158));
DFF_X1 \Acc_reg[9]  (.Q (\Acc[9] ), .CK (CTS_n_tid0_49), .D (n_159));
DFF_X1 \Acc_reg[10]  (.Q (\Acc[10] ), .CK (CTS_n_tid0_49), .D (n_160));
DFF_X1 \Acc_reg[11]  (.Q (\Acc[11] ), .CK (CTS_n_tid0_49), .D (n_161));
DFF_X1 \Acc_reg[12]  (.Q (\Acc[12] ), .CK (CTS_n_tid0_49), .D (n_162));
DFF_X1 \Acc_reg[13]  (.Q (\Acc[13] ), .CK (CTS_n_tid0_49), .D (n_163));
DFF_X1 \Acc_reg[14]  (.Q (\Acc[14] ), .CK (CTS_n_tid0_49), .D (n_164));
DFF_X1 \Acc_reg[15]  (.Q (\Acc[15] ), .CK (CTS_n_tid0_49), .D (n_165));
DFF_X1 \Acc_reg[16]  (.Q (\Acc[16] ), .CK (CTS_n_tid0_49), .D (n_166));
DFF_X1 \Acc_reg[17]  (.Q (\Acc[17] ), .CK (CTS_n_tid0_49), .D (n_168));
DFF_X1 \Acc_reg[18]  (.Q (\Acc[18] ), .CK (CTS_n_tid0_49), .D (n_169));
DFF_X1 \Acc_reg[19]  (.Q (\Acc[19] ), .CK (CTS_n_tid0_49), .D (n_170));
DFF_X1 \Acc_reg[20]  (.Q (\Acc[20] ), .CK (CTS_n_tid0_49), .D (n_171));
DFF_X1 \Acc_reg[21]  (.Q (\Acc[21] ), .CK (CTS_n_tid0_49), .D (n_172));
DFF_X1 \Acc_reg[22]  (.Q (\Acc[22] ), .CK (CTS_n_tid0_49), .D (n_173));
DFF_X1 \Acc_reg[23]  (.Q (\Acc[23] ), .CK (CTS_n_tid0_49), .D (n_174));
DFF_X1 \Acc_reg[24]  (.Q (\Acc[24] ), .CK (CTS_n_tid0_49), .D (n_175));
DFF_X1 \Acc_reg[25]  (.Q (\Acc[25] ), .CK (CTS_n_tid0_49), .D (n_176));
DFF_X1 \Acc_reg[26]  (.Q (\Acc[26] ), .CK (CTS_n_tid0_49), .D (n_177));
DFF_X1 \Acc_reg[27]  (.Q (\Acc[27] ), .CK (CTS_n_tid0_49), .D (n_178));
DFF_X1 \Acc_reg[28]  (.Q (\Acc[28] ), .CK (CTS_n_tid0_49), .D (n_179));
DFF_X1 \Acc_reg[29]  (.Q (\Acc[29] ), .CK (CTS_n_tid0_49), .D (n_180));
DFF_X1 \Acc_reg[30]  (.Q (\Acc[30] ), .CK (CTS_n_tid0_49), .D (n_181));
DFF_X1 \Acc_reg[31]  (.Q (\Acc[31] ), .CK (CTS_n_tid0_49), .D (n_182));
CLKGATETST_X8 clk_gate_Acc_reg (.GCK (CTS_n_tid0_56), .CK (CTS_n_tid0_209), .E (n_149), .SE (1'b0 ));
DFF_X1 \inputQ_reg_reg[0]  (.Q (\inputQ_reg[0] ), .CK (n_133), .D (n_184));
DFF_X1 \inputQ_reg_reg[1]  (.Q (\inputQ_reg[1] ), .CK (n_133), .D (n_185));
DFF_X1 \inputQ_reg_reg[2]  (.Q (\inputQ_reg[2] ), .CK (n_133), .D (n_186));
DFF_X1 \inputQ_reg_reg[3]  (.Q (\inputQ_reg[3] ), .CK (n_133), .D (n_187));
DFF_X1 \inputQ_reg_reg[4]  (.Q (\inputQ_reg[4] ), .CK (n_133), .D (n_188));
DFF_X1 \inputQ_reg_reg[5]  (.Q (\inputQ_reg[5] ), .CK (n_133), .D (n_189));
DFF_X1 \inputQ_reg_reg[6]  (.Q (\inputQ_reg[6] ), .CK (n_133), .D (n_190));
DFF_X1 \inputQ_reg_reg[7]  (.Q (\inputQ_reg[7] ), .CK (n_133), .D (n_191));
DFF_X1 \inputQ_reg_reg[8]  (.Q (\inputQ_reg[8] ), .CK (n_133), .D (n_192));
DFF_X1 \inputQ_reg_reg[9]  (.Q (\inputQ_reg[9] ), .CK (n_133), .D (n_193));
DFF_X1 \inputQ_reg_reg[10]  (.Q (\inputQ_reg[10] ), .CK (n_133), .D (n_194));
DFF_X1 \inputQ_reg_reg[11]  (.Q (\inputQ_reg[11] ), .CK (n_133), .D (n_195));
DFF_X1 \inputQ_reg_reg[12]  (.Q (\inputQ_reg[12] ), .CK (n_133), .D (n_196));
DFF_X1 \inputQ_reg_reg[13]  (.Q (\inputQ_reg[13] ), .CK (n_133), .D (n_197));
DFF_X1 \inputQ_reg_reg[14]  (.Q (\inputQ_reg[14] ), .CK (n_133), .D (n_198));
DFF_X1 \inputQ_reg_reg[15]  (.Q (\inputQ_reg[15] ), .CK (n_133), .D (n_199));
DFF_X1 \inputQ_reg_reg[16]  (.Q (\inputQ_reg[16] ), .CK (n_133), .D (n_200));
DFF_X1 \inputQ_reg_reg[17]  (.Q (\inputQ_reg[17] ), .CK (n_133), .D (n_202));
DFF_X1 \inputQ_reg_reg[18]  (.Q (\inputQ_reg[18] ), .CK (n_133), .D (n_203));
DFF_X1 \inputQ_reg_reg[19]  (.Q (\inputQ_reg[19] ), .CK (n_133), .D (n_204));
DFF_X1 \inputQ_reg_reg[20]  (.Q (\inputQ_reg[20] ), .CK (n_133), .D (n_205));
DFF_X1 \inputQ_reg_reg[21]  (.Q (\inputQ_reg[21] ), .CK (n_133), .D (n_206));
DFF_X1 \inputQ_reg_reg[22]  (.Q (\inputQ_reg[22] ), .CK (n_133), .D (n_207));
DFF_X1 \inputQ_reg_reg[23]  (.Q (\inputQ_reg[23] ), .CK (n_133), .D (n_208));
DFF_X1 \inputQ_reg_reg[24]  (.Q (\inputQ_reg[24] ), .CK (n_133), .D (n_209));
DFF_X1 \inputQ_reg_reg[25]  (.Q (\inputQ_reg[25] ), .CK (n_133), .D (n_210));
DFF_X1 \inputQ_reg_reg[26]  (.Q (\inputQ_reg[26] ), .CK (n_133), .D (n_211));
DFF_X1 \inputQ_reg_reg[27]  (.Q (\inputQ_reg[27] ), .CK (n_133), .D (n_212));
DFF_X1 \inputQ_reg_reg[28]  (.Q (\inputQ_reg[28] ), .CK (n_133), .D (n_213));
DFF_X1 \inputQ_reg_reg[29]  (.Q (\inputQ_reg[29] ), .CK (n_133), .D (n_214));
DFF_X1 \inputQ_reg_reg[30]  (.Q (\inputQ_reg[30] ), .CK (n_133), .D (n_215));
DFF_X1 \inputQ_reg_reg[31]  (.Q (\inputQ_reg[31] ), .CK (n_133), .D (n_216));
CLKGATETST_X1 clk_gate_inputQ_reg_reg (.GCK (n_133), .CK (clk_CTS_0_PP_0), .E (n_183), .SE (1'b0 ));
datapath i_0 (.p_0 ({n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
    n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
    n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, 
    n_2}), .input_plus (input_plus), .p_1 ({\Acc[31] , \Acc[30] , \Acc[29] , \Acc[28] , 
    \Acc[27] , \Acc[26] , \Acc[25] , \Acc[24] , \Acc[23] , \Acc[22] , \Acc[21] , 
    \Acc[20] , \Acc[19] , \Acc[18] , \Acc[17] , \Acc[16] , \Acc[15] , \Acc[14] , 
    \Acc[13] , \Acc[12] , \Acc[11] , \Acc[10] , \Acc[9] , \Acc[8] , \Acc[7] , \Acc[6] , 
    \Acc[5] , \Acc[4] , \Acc[3] , \Acc[2] , \Acc[1] , \Acc[0] , \inputQ_reg[31] , 
    \inputQ_reg[30] , \inputQ_reg[29] , \inputQ_reg[28] , \inputQ_reg[27] , \inputQ_reg[26] , 
    \inputQ_reg[25] , \inputQ_reg[24] , \inputQ_reg[23] , \inputQ_reg[22] , \inputQ_reg[21] , 
    \inputQ_reg[20] , \inputQ_reg[19] , \inputQ_reg[18] , \inputQ_reg[17] , \inputQ_reg[16] , 
    \inputQ_reg[15] , \inputQ_reg[14] , \inputQ_reg[13] , \inputQ_reg[12] , \inputQ_reg[11] , 
    \inputQ_reg[10] , \inputQ_reg[9] , \inputQ_reg[8] , \inputQ_reg[7] , \inputQ_reg[6] , 
    \inputQ_reg[5] , \inputQ_reg[4] , \inputQ_reg[3] , \inputQ_reg[2] , \inputQ_reg[1] , 
    \inputQ_reg[0] }));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_121), .D (n_219));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_121), .D (n_220));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_121), .D (n_221));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid0_121), .D (n_222));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid0_121), .D (n_223));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid0_121), .D (n_224));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_121), .D (n_225));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid0_121), .D (n_226));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid0_121), .D (n_227));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid0_121), .D (n_228));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid0_121), .D (n_229));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid0_121), .D (n_230));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid0_121), .D (n_231));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_121), .D (n_232));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_121), .D (n_233));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_121), .D (n_234));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_121), .D (n_235));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_122), .D (n_236));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_122), .D (n_237));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_122), .D (n_238));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_122), .D (n_239));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_122), .D (n_240));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_122), .D (n_241));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_122), .D (n_242));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_122), .D (n_243));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_122), .D (n_244));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_122), .D (n_245));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_122), .D (n_246));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_122), .D (n_247));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_122), .D (n_248));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_122), .D (n_249));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid0_122), .D (n_250));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n_tid0_122), .D (n_251));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n_tid0_122), .D (n_252));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n_tid0_122), .D (n_253));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n_tid0_122), .D (n_254));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n_tid0_122), .D (n_255));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n_tid0_122), .D (n_256));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n_tid0_112), .D (n_257));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n_tid0_112), .D (n_258));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n_tid0_112), .D (n_259));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n_tid0_112), .D (n_260));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n_tid0_112), .D (n_261));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n_tid0_112), .D (n_262));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n_tid0_112), .D (n_263));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n_tid0_112), .D (n_264));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n_tid0_112), .D (n_265));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n_tid0_112), .D (n_266));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n_tid0_112), .D (n_267));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n_tid0_112), .D (n_268));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n_tid0_112), .D (n_269));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n_tid0_112), .D (n_270));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n_tid0_112), .D (n_271));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n_tid0_112), .D (n_272));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n_tid0_112), .D (n_273));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n_tid0_112), .D (n_274));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n_tid0_112), .D (n_275));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n_tid0_112), .D (n_276));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n_tid0_112), .D (n_277));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n_tid0_112), .D (n_278));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n_tid0_112), .D (n_279));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n_tid0_112), .D (n_280));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (CTS_n_tid0_112), .D (n_281));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n_tid0_112), .D (n_282));
CLKBUF_X2 hfn_ipo_c9 (.Z (hfn_ipo_n9), .A (n_2_115));
CLKBUF_X2 hfn_ipo_c10 (.Z (hfn_ipo_n10), .A (n_2_115));
CLKBUF_X2 hfn_ipo_c11 (.Z (hfn_ipo_n11), .A (n_2_116));
CLKBUF_X2 hfn_ipo_c12 (.Z (hfn_ipo_n12), .A (n_2_116));
CLKBUF_X3 CTS_L4_c_tid1_23 (.Z (CTS_n_tid1_16), .A (CTS_n_tid1_17));
CLKBUF_X3 CTS_L4_c_tid0_85 (.Z (CTS_n_tid0_112), .A (CTS_n_tid0_188));
CLKBUF_X1 CTS_L2_c_tid0_164 (.Z (CTS_n_tid0_209), .A (clk_CTS_0_PP_0));
CLKBUF_X3 CTS_L4_c_tid0_39 (.Z (CTS_n_tid0_49), .A (CTS_n_tid0_56));
CLKBUF_X2 CTS_L4_c_tid0_94 (.Z (CTS_n_tid0_121), .A (CTS_n_tid0_188));
CLKBUF_X2 CTS_L4_c_tid0_95 (.Z (CTS_n_tid0_122), .A (CTS_n_tid0_188));
CLKBUF_X1 CTS_L1_c_tid0_175 (.Z (clk_CTS_0_PP_0), .A (clk_CTS_0_PP_1));
CLKBUF_X1 CTS_L3_c_tid0_153 (.Z (CTS_n_tid0_198), .A (CTS_n_tid0_209));

endmodule //controller

module multiplier (clk, reset, en, inputM, inputQ, input_plus, out);

output [63:0] out;
input clk;
input en;
input [31:0] inputM;
input [31:0] inputQ;
input input_plus;
input reset;
wire CTS_n_tid0_3;
wire \preout[63] ;
wire \preout[62] ;
wire \preout[61] ;
wire \preout[60] ;
wire \preout[59] ;
wire \preout[58] ;
wire \preout[57] ;
wire \preout[56] ;
wire \preout[55] ;
wire \preout[54] ;
wire \preout[53] ;
wire \preout[52] ;
wire \preout[51] ;
wire \preout[50] ;
wire \preout[49] ;
wire \preout[48] ;
wire \preout[47] ;
wire \preout[46] ;
wire \preout[45] ;
wire \preout[44] ;
wire \preout[43] ;
wire \preout[42] ;
wire \preout[41] ;
wire \preout[40] ;
wire \preout[39] ;
wire \preout[38] ;
wire \preout[37] ;
wire \preout[36] ;
wire \preout[35] ;
wire \preout[34] ;
wire \preout[33] ;
wire \preout[32] ;
wire \preout[31] ;
wire \preout[30] ;
wire \preout[29] ;
wire \preout[28] ;
wire \preout[27] ;
wire \preout[26] ;
wire \preout[25] ;
wire \preout[24] ;
wire \preout[23] ;
wire \preout[22] ;
wire \preout[21] ;
wire \preout[20] ;
wire \preout[19] ;
wire \preout[18] ;
wire \preout[17] ;
wire \preout[16] ;
wire \preout[15] ;
wire \preout[14] ;
wire \preout[13] ;
wire \preout[12] ;
wire \preout[11] ;
wire \preout[10] ;
wire \preout[9] ;
wire \preout[8] ;
wire \preout[7] ;
wire \preout[6] ;
wire \preout[5] ;
wire \preout[4] ;
wire \preout[3] ;
wire \preout[2] ;
wire \preout[1] ;
wire \preout[0] ;
wire \inputQ_inv22[31] ;
wire \inputQ_inv22[30] ;
wire \inputQ_inv22[29] ;
wire \inputQ_inv22[28] ;
wire \inputQ_inv22[27] ;
wire \inputQ_inv22[26] ;
wire \inputQ_inv22[25] ;
wire \inputQ_inv22[24] ;
wire \inputQ_inv22[23] ;
wire \inputQ_inv22[22] ;
wire \inputQ_inv22[21] ;
wire \inputQ_inv22[20] ;
wire \inputQ_inv22[19] ;
wire \inputQ_inv22[18] ;
wire \inputQ_inv22[17] ;
wire \inputQ_inv22[16] ;
wire \inputQ_inv22[15] ;
wire \inputQ_inv22[14] ;
wire \inputQ_inv22[13] ;
wire \inputQ_inv22[12] ;
wire \inputQ_inv22[11] ;
wire \inputQ_inv22[10] ;
wire \inputQ_inv22[9] ;
wire \inputQ_inv22[8] ;
wire \inputQ_inv22[7] ;
wire \inputQ_inv22[6] ;
wire \inputQ_inv22[5] ;
wire \inputQ_inv22[4] ;
wire \inputQ_inv22[3] ;
wire \inputQ_inv22[2] ;
wire \inputQ_inv22[1] ;
wire \inputQ_inv22[0] ;
wire \inputM_inv22[31] ;
wire \inputM_inv22[30] ;
wire \inputM_inv22[29] ;
wire \inputM_inv22[28] ;
wire \inputM_inv22[27] ;
wire \inputM_inv22[26] ;
wire \inputM_inv22[25] ;
wire \inputM_inv22[24] ;
wire \inputM_inv22[23] ;
wire \inputM_inv22[22] ;
wire \inputM_inv22[21] ;
wire \inputM_inv22[20] ;
wire \inputM_inv22[19] ;
wire \inputM_inv22[18] ;
wire \inputM_inv22[17] ;
wire \inputM_inv22[16] ;
wire \inputM_inv22[15] ;
wire \inputM_inv22[14] ;
wire \inputM_inv22[13] ;
wire \inputM_inv22[12] ;
wire \inputM_inv22[11] ;
wire \inputM_inv22[10] ;
wire \inputM_inv22[9] ;
wire \inputM_inv22[8] ;
wire \inputM_inv22[7] ;
wire \inputM_inv22[6] ;
wire \inputM_inv22[5] ;
wire \inputM_inv22[4] ;
wire \inputM_inv22[3] ;
wire \inputM_inv22[2] ;
wire \inputM_inv22[1] ;
wire \inputM_inv22[0] ;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;


AND2_X1 i_0_1_63 (.ZN (n_0_63), .A1 (\inputM_inv22[31] ), .A2 (inputM[31]));
MUX2_X1 i_0_1_62 (.Z (n_0_62), .A (inputM[30]), .B (\inputM_inv22[30] ), .S (inputM[31]));
MUX2_X1 i_0_1_61 (.Z (n_0_61), .A (inputM[29]), .B (\inputM_inv22[29] ), .S (inputM[31]));
MUX2_X1 i_0_1_60 (.Z (n_0_60), .A (inputM[28]), .B (\inputM_inv22[28] ), .S (inputM[31]));
MUX2_X1 i_0_1_59 (.Z (n_0_59), .A (inputM[27]), .B (\inputM_inv22[27] ), .S (inputM[31]));
MUX2_X1 i_0_1_58 (.Z (n_0_58), .A (inputM[26]), .B (\inputM_inv22[26] ), .S (inputM[31]));
MUX2_X1 i_0_1_57 (.Z (n_0_57), .A (inputM[25]), .B (\inputM_inv22[25] ), .S (inputM[31]));
MUX2_X1 i_0_1_56 (.Z (n_0_56), .A (inputM[24]), .B (\inputM_inv22[24] ), .S (inputM[31]));
MUX2_X1 i_0_1_55 (.Z (n_0_55), .A (inputM[23]), .B (\inputM_inv22[23] ), .S (inputM[31]));
MUX2_X1 i_0_1_54 (.Z (n_0_54), .A (inputM[22]), .B (\inputM_inv22[22] ), .S (inputM[31]));
MUX2_X1 i_0_1_53 (.Z (n_0_53), .A (inputM[21]), .B (\inputM_inv22[21] ), .S (inputM[31]));
MUX2_X1 i_0_1_52 (.Z (n_0_52), .A (inputM[20]), .B (\inputM_inv22[20] ), .S (inputM[31]));
MUX2_X1 i_0_1_51 (.Z (n_0_51), .A (inputM[19]), .B (\inputM_inv22[19] ), .S (inputM[31]));
MUX2_X1 i_0_1_50 (.Z (n_0_50), .A (inputM[18]), .B (\inputM_inv22[18] ), .S (inputM[31]));
MUX2_X1 i_0_1_49 (.Z (n_0_49), .A (inputM[17]), .B (\inputM_inv22[17] ), .S (inputM[31]));
MUX2_X1 i_0_1_48 (.Z (n_0_48), .A (inputM[16]), .B (\inputM_inv22[16] ), .S (inputM[31]));
MUX2_X1 i_0_1_47 (.Z (n_0_47), .A (inputM[15]), .B (\inputM_inv22[15] ), .S (inputM[31]));
MUX2_X1 i_0_1_46 (.Z (n_0_46), .A (inputM[14]), .B (\inputM_inv22[14] ), .S (inputM[31]));
MUX2_X1 i_0_1_45 (.Z (n_0_45), .A (inputM[13]), .B (\inputM_inv22[13] ), .S (inputM[31]));
MUX2_X1 i_0_1_44 (.Z (n_0_44), .A (inputM[12]), .B (\inputM_inv22[12] ), .S (inputM[31]));
MUX2_X1 i_0_1_43 (.Z (n_0_43), .A (inputM[11]), .B (\inputM_inv22[11] ), .S (inputM[31]));
MUX2_X1 i_0_1_42 (.Z (n_0_42), .A (inputM[10]), .B (\inputM_inv22[10] ), .S (inputM[31]));
MUX2_X1 i_0_1_41 (.Z (n_0_41), .A (inputM[9]), .B (\inputM_inv22[9] ), .S (inputM[31]));
MUX2_X1 i_0_1_40 (.Z (n_0_40), .A (inputM[8]), .B (\inputM_inv22[8] ), .S (inputM[31]));
MUX2_X1 i_0_1_39 (.Z (n_0_39), .A (inputM[7]), .B (\inputM_inv22[7] ), .S (inputM[31]));
MUX2_X1 i_0_1_38 (.Z (n_0_38), .A (inputM[6]), .B (\inputM_inv22[6] ), .S (inputM[31]));
MUX2_X1 i_0_1_37 (.Z (n_0_37), .A (inputM[5]), .B (\inputM_inv22[5] ), .S (inputM[31]));
MUX2_X1 i_0_1_36 (.Z (n_0_36), .A (inputM[4]), .B (\inputM_inv22[4] ), .S (inputM[31]));
MUX2_X1 i_0_1_35 (.Z (n_0_35), .A (inputM[3]), .B (\inputM_inv22[3] ), .S (inputM[31]));
MUX2_X1 i_0_1_34 (.Z (n_0_34), .A (inputM[2]), .B (\inputM_inv22[2] ), .S (inputM[31]));
MUX2_X1 i_0_1_33 (.Z (n_0_33), .A (inputM[1]), .B (\inputM_inv22[1] ), .S (inputM[31]));
MUX2_X1 i_0_1_32 (.Z (n_0_32), .A (inputM[0]), .B (\inputM_inv22[0] ), .S (inputM[31]));
AND2_X1 i_0_1_31 (.ZN (n_0_31), .A1 (\inputQ_inv22[31] ), .A2 (inputQ[31]));
MUX2_X1 i_0_1_30 (.Z (n_0_30), .A (inputQ[30]), .B (\inputQ_inv22[30] ), .S (inputQ[31]));
MUX2_X1 i_0_1_29 (.Z (n_0_29), .A (inputQ[29]), .B (\inputQ_inv22[29] ), .S (inputQ[31]));
MUX2_X1 i_0_1_28 (.Z (n_0_28), .A (inputQ[28]), .B (\inputQ_inv22[28] ), .S (inputQ[31]));
MUX2_X1 i_0_1_27 (.Z (n_0_27), .A (inputQ[27]), .B (\inputQ_inv22[27] ), .S (inputQ[31]));
MUX2_X1 i_0_1_26 (.Z (n_0_26), .A (inputQ[26]), .B (\inputQ_inv22[26] ), .S (inputQ[31]));
MUX2_X1 i_0_1_25 (.Z (n_0_25), .A (inputQ[25]), .B (\inputQ_inv22[25] ), .S (inputQ[31]));
MUX2_X1 i_0_1_24 (.Z (n_0_24), .A (inputQ[24]), .B (\inputQ_inv22[24] ), .S (inputQ[31]));
MUX2_X1 i_0_1_23 (.Z (n_0_23), .A (inputQ[23]), .B (\inputQ_inv22[23] ), .S (inputQ[31]));
MUX2_X1 i_0_1_22 (.Z (n_0_22), .A (inputQ[22]), .B (\inputQ_inv22[22] ), .S (inputQ[31]));
MUX2_X1 i_0_1_21 (.Z (n_0_21), .A (inputQ[21]), .B (\inputQ_inv22[21] ), .S (inputQ[31]));
MUX2_X1 i_0_1_20 (.Z (n_0_20), .A (inputQ[20]), .B (\inputQ_inv22[20] ), .S (inputQ[31]));
MUX2_X1 i_0_1_19 (.Z (n_0_19), .A (inputQ[19]), .B (\inputQ_inv22[19] ), .S (inputQ[31]));
MUX2_X1 i_0_1_18 (.Z (n_0_18), .A (inputQ[18]), .B (\inputQ_inv22[18] ), .S (inputQ[31]));
MUX2_X1 i_0_1_17 (.Z (n_0_17), .A (inputQ[17]), .B (\inputQ_inv22[17] ), .S (inputQ[31]));
MUX2_X1 i_0_1_16 (.Z (n_0_16), .A (inputQ[16]), .B (\inputQ_inv22[16] ), .S (inputQ[31]));
MUX2_X1 i_0_1_15 (.Z (n_0_15), .A (inputQ[15]), .B (\inputQ_inv22[15] ), .S (inputQ[31]));
MUX2_X1 i_0_1_14 (.Z (n_0_14), .A (inputQ[14]), .B (\inputQ_inv22[14] ), .S (inputQ[31]));
MUX2_X1 i_0_1_13 (.Z (n_0_13), .A (inputQ[13]), .B (\inputQ_inv22[13] ), .S (inputQ[31]));
MUX2_X1 i_0_1_12 (.Z (n_0_12), .A (inputQ[12]), .B (\inputQ_inv22[12] ), .S (inputQ[31]));
MUX2_X1 i_0_1_11 (.Z (n_0_11), .A (inputQ[11]), .B (\inputQ_inv22[11] ), .S (inputQ[31]));
MUX2_X1 i_0_1_10 (.Z (n_0_10), .A (inputQ[10]), .B (\inputQ_inv22[10] ), .S (inputQ[31]));
MUX2_X1 i_0_1_9 (.Z (n_0_9), .A (inputQ[9]), .B (\inputQ_inv22[9] ), .S (inputQ[31]));
MUX2_X1 i_0_1_8 (.Z (n_0_8), .A (inputQ[8]), .B (\inputQ_inv22[8] ), .S (inputQ[31]));
MUX2_X1 i_0_1_7 (.Z (n_0_7), .A (inputQ[7]), .B (\inputQ_inv22[7] ), .S (inputQ[31]));
MUX2_X1 i_0_1_6 (.Z (n_0_6), .A (inputQ[6]), .B (\inputQ_inv22[6] ), .S (inputQ[31]));
MUX2_X1 i_0_1_5 (.Z (n_0_5), .A (inputQ[5]), .B (\inputQ_inv22[5] ), .S (inputQ[31]));
MUX2_X1 i_0_1_4 (.Z (n_0_4), .A (inputQ[4]), .B (\inputQ_inv22[4] ), .S (inputQ[31]));
MUX2_X1 i_0_1_3 (.Z (n_0_3), .A (inputQ[3]), .B (\inputQ_inv22[3] ), .S (inputQ[31]));
MUX2_X1 i_0_1_2 (.Z (n_0_2), .A (inputQ[2]), .B (\inputQ_inv22[2] ), .S (inputQ[31]));
MUX2_X1 i_0_1_1 (.Z (n_0_1), .A (inputQ[1]), .B (\inputQ_inv22[1] ), .S (inputQ[31]));
MUX2_X1 i_0_1_0 (.Z (n_0_0), .A (inputQ[0]), .B (\inputQ_inv22[0] ), .S (inputQ[31]));
datapath__0_29 i_0_2 (.inputM_inv22 ({\inputM_inv22[31] , \inputM_inv22[30] , \inputM_inv22[29] , 
    \inputM_inv22[28] , \inputM_inv22[27] , \inputM_inv22[26] , \inputM_inv22[25] , 
    \inputM_inv22[24] , \inputM_inv22[23] , \inputM_inv22[22] , \inputM_inv22[21] , 
    \inputM_inv22[20] , \inputM_inv22[19] , \inputM_inv22[18] , \inputM_inv22[17] , 
    \inputM_inv22[16] , \inputM_inv22[15] , \inputM_inv22[14] , \inputM_inv22[13] , 
    \inputM_inv22[12] , \inputM_inv22[11] , \inputM_inv22[10] , \inputM_inv22[9] , 
    \inputM_inv22[8] , \inputM_inv22[7] , \inputM_inv22[6] , \inputM_inv22[5] , \inputM_inv22[4] , 
    \inputM_inv22[3] , \inputM_inv22[2] , \inputM_inv22[1] , \inputM_inv22[0] }), .inputM ({
    inputM[31], inputM[30], inputM[29], inputM[28], inputM[27], inputM[26], inputM[25], 
    inputM[24], inputM[23], inputM[22], inputM[21], inputM[20], inputM[19], inputM[18], 
    inputM[17], inputM[16], inputM[15], inputM[14], inputM[13], inputM[12], inputM[11], 
    inputM[10], inputM[9], inputM[8], inputM[7], inputM[6], inputM[5], inputM[4], 
    inputM[3], inputM[2], inputM[1], inputM[0]}), .input_plus (input_plus));
datapath__0_27 i_0_0 (.inputQ_inv22 ({\inputQ_inv22[31] , \inputQ_inv22[30] , \inputQ_inv22[29] , 
    \inputQ_inv22[28] , \inputQ_inv22[27] , \inputQ_inv22[26] , \inputQ_inv22[25] , 
    \inputQ_inv22[24] , \inputQ_inv22[23] , \inputQ_inv22[22] , \inputQ_inv22[21] , 
    \inputQ_inv22[20] , \inputQ_inv22[19] , \inputQ_inv22[18] , \inputQ_inv22[17] , 
    \inputQ_inv22[16] , \inputQ_inv22[15] , \inputQ_inv22[14] , \inputQ_inv22[13] , 
    \inputQ_inv22[12] , \inputQ_inv22[11] , \inputQ_inv22[10] , \inputQ_inv22[9] , 
    \inputQ_inv22[8] , \inputQ_inv22[7] , \inputQ_inv22[6] , \inputQ_inv22[5] , \inputQ_inv22[4] , 
    \inputQ_inv22[3] , \inputQ_inv22[2] , \inputQ_inv22[1] , \inputQ_inv22[0] }), .inputQ ({
    inputQ[31], inputQ[30], inputQ[29], inputQ[28], inputQ[27], inputQ[26], inputQ[25], 
    inputQ[24], inputQ[23], inputQ[22], inputQ[21], inputQ[20], inputQ[19], inputQ[18], 
    inputQ[17], inputQ[16], inputQ[15], inputQ[14], inputQ[13], inputQ[12], inputQ[11], 
    inputQ[10], inputQ[9], inputQ[8], inputQ[7], inputQ[6], inputQ[5], inputQ[4], 
    inputQ[3], inputQ[2], inputQ[1], inputQ[0]}), .input_plus (input_plus));
registerNbits__parameterized0 reg3 (.out ({out[63], out[62], out[61], out[60], out[59], 
    out[58], out[57], out[56], out[55], out[54], out[53], out[52], out[51], out[50], 
    out[49], out[48], out[47], out[46], out[45], out[44], out[43], out[42], out[41], 
    out[40], out[39], out[38], out[37], out[36], out[35], out[34], out[33], out[32], 
    out[31], out[30], out[29], out[28], out[27], out[26], out[25], out[24], out[23], 
    out[22], out[21], out[20], out[19], out[18], out[17], out[16], out[15], out[14], 
    out[13], out[12], out[11], out[10], out[9], out[8], out[7], out[6], out[5], out[4], 
    out[3], out[2], out[1], out[0]}), .en (en), .inp ({\preout[63] , \preout[62] , 
    \preout[61] , \preout[60] , \preout[59] , \preout[58] , \preout[57] , \preout[56] , 
    \preout[55] , \preout[54] , \preout[53] , \preout[52] , \preout[51] , \preout[50] , 
    \preout[49] , \preout[48] , \preout[47] , \preout[46] , \preout[45] , \preout[44] , 
    \preout[43] , \preout[42] , \preout[41] , \preout[40] , \preout[39] , \preout[38] , 
    \preout[37] , \preout[36] , \preout[35] , \preout[34] , \preout[33] , \preout[32] , 
    \preout[31] , \preout[30] , \preout[29] , \preout[28] , \preout[27] , \preout[26] , 
    \preout[25] , \preout[24] , \preout[23] , \preout[22] , \preout[21] , \preout[20] , 
    \preout[19] , \preout[18] , \preout[17] , \preout[16] , \preout[15] , \preout[14] , 
    \preout[13] , \preout[12] , \preout[11] , \preout[10] , \preout[9] , \preout[8] , 
    \preout[7] , \preout[6] , \preout[5] , \preout[4] , \preout[3] , \preout[2] , 
    \preout[1] , \preout[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_3));
controller controller (.out ({\preout[63] , \preout[62] , \preout[61] , \preout[60] , 
    \preout[59] , \preout[58] , \preout[57] , \preout[56] , \preout[55] , \preout[54] , 
    \preout[53] , \preout[52] , \preout[51] , \preout[50] , \preout[49] , \preout[48] , 
    \preout[47] , \preout[46] , \preout[45] , \preout[44] , \preout[43] , \preout[42] , 
    \preout[41] , \preout[40] , \preout[39] , \preout[38] , \preout[37] , \preout[36] , 
    \preout[35] , \preout[34] , \preout[33] , \preout[32] , \preout[31] , \preout[30] , 
    \preout[29] , \preout[28] , \preout[27] , \preout[26] , \preout[25] , \preout[24] , 
    \preout[23] , \preout[22] , \preout[21] , \preout[20] , \preout[19] , \preout[18] , 
    \preout[17] , \preout[16] , \preout[15] , \preout[14] , \preout[13] , \preout[12] , 
    \preout[11] , \preout[10] , \preout[9] , \preout[8] , \preout[7] , \preout[6] , 
    \preout[5] , \preout[4] , \preout[3] , \preout[2] , \preout[1] , \preout[0] })
    , .clk_CTS_0_PP_0 (CTS_n_tid0_3), .Mbit (inputM[31]), .Qbit (inputQ[31]), .inputM_wire ({
    n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
    n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, 
    n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, 
    n_0_33, n_0_32}), .inputQ_wire ({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
    n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
    n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
    n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}), .input_plus (input_plus), .reset (reset)
    , .clk_CTS_0_PP_1 (clk));

endmodule //multiplier


