
// 	Sat Dec 24 10:29:18 2022
//	vlsi
//	localhost.localdomain

module datapath__0_195 (p_0, p_1);

output [32:0] p_0;
input [32:0] p_1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (p_1[25]));
INV_X1 i_63 (.ZN (n_32), .A (p_1[21]));
INV_X1 i_62 (.ZN (n_31), .A (p_1[14]));
INV_X1 i_61 (.ZN (n_30), .A (p_1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (p_1[2]), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (p_1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (p_1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (p_1[5]), .A3 (p_1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (p_1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (p_1[8]), .A3 (p_1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (p_1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (p_1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (p_1[12]), .A3 (p_1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (p_1[15]), .A3 (p_1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (p_1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (p_1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]), .A4 (p_1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (p_1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (p_1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (p_1[23]), .A3 (p_1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (p_1[26]), .A3 (p_1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (p_1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]), .A4 (p_1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (p_1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (p_1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (p_1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (p_1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (p_1[27]), .B1 (n_9), .B2 (p_1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (p_1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (p_1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (p_1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (p_1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (p_1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (p_1[16]), .B1 (n_19), .B2 (p_1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (p_1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (p_1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (p_1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (p_1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (p_1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (p_1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[9]), .B1 (n_25), .B2 (p_1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (p_1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (p_1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[6]), .B1 (n_27), .B2 (p_1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (p_1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (p_1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (p_1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[2]), .B1 (p_1[1]), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (p_1[1]), .B (p_1[0]));

endmodule //datapath__0_195

module datapath__0_193 (p_0, read_data2);

output [31:0] p_0;
input [31:0] read_data2;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (read_data2[25]));
INV_X1 i_63 (.ZN (n_32), .A (read_data2[21]));
INV_X1 i_62 (.ZN (n_31), .A (read_data2[14]));
INV_X1 i_61 (.ZN (n_30), .A (read_data2[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (read_data2[2]), .A2 (read_data2[1]), .A3 (read_data2[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (read_data2[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (read_data2[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (read_data2[5]), .A3 (read_data2[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (read_data2[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (read_data2[8]), .A3 (read_data2[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (read_data2[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (read_data2[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (read_data2[12]), .A3 (read_data2[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (read_data2[15]), .A3 (read_data2[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (read_data2[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (read_data2[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (read_data2[18]), .A3 (read_data2[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (read_data2[18]), .A3 (read_data2[19]), .A4 (read_data2[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (read_data2[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (read_data2[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (read_data2[23]), .A3 (read_data2[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (read_data2[26]), .A3 (read_data2[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (read_data2[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (read_data2[28]), .A3 (read_data2[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (read_data2[28]), .A3 (read_data2[29]), .A4 (read_data2[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (read_data2[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (read_data2[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (read_data2[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (read_data2[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (read_data2[27]), .B1 (n_9), .B2 (read_data2[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (read_data2[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (read_data2[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (read_data2[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (read_data2[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (read_data2[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (read_data2[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (read_data2[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (read_data2[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (read_data2[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (read_data2[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (read_data2[16]), .B1 (n_19), .B2 (read_data2[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (read_data2[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (read_data2[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (read_data2[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (read_data2[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (read_data2[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (read_data2[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (read_data2[9]), .B1 (n_25), .B2 (read_data2[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (read_data2[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (read_data2[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (read_data2[6]), .B1 (n_27), .B2 (read_data2[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (read_data2[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (read_data2[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (read_data2[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (read_data2[2]), .B1 (read_data2[1]), .B2 (read_data2[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (read_data2[1]), .B (read_data2[0]));

endmodule //datapath__0_193

module regFile64 (clk__CTS_1_PP_1, read_data, write_en, write_data, clk);

output [63:0] read_data;
input clk;
input [63:0] write_data;
input write_en;
input clk__CTS_1_PP_1;
wire CTS_n_tid1_7;
wire n_tid1_34;


DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid1_7), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid1_7), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid1_7), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid1_7), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid1_7), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid1_7), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid1_7), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid1_7), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid1_7), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid1_7), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid1_7), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid1_7), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid1_7), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid1_7), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid1_7), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid1_7), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid1_7), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid1_7), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid1_7), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid1_7), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid1_7), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid1_7), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid1_7), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid1_7), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid1_7), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid1_7), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid1_7), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid1_7), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid1_7), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid1_7), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid1_7), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid1_7), .D (write_data[31]));
DFF_X1 \my_reg_reg[32]  (.Q (read_data[32]), .CK (CTS_n_tid1_7), .D (write_data[32]));
DFF_X1 \my_reg_reg[33]  (.Q (read_data[33]), .CK (CTS_n_tid1_7), .D (write_data[33]));
DFF_X1 \my_reg_reg[34]  (.Q (read_data[34]), .CK (CTS_n_tid1_7), .D (write_data[34]));
DFF_X1 \my_reg_reg[35]  (.Q (read_data[35]), .CK (CTS_n_tid1_7), .D (write_data[35]));
DFF_X1 \my_reg_reg[36]  (.Q (read_data[36]), .CK (CTS_n_tid1_7), .D (write_data[36]));
DFF_X1 \my_reg_reg[37]  (.Q (read_data[37]), .CK (CTS_n_tid1_7), .D (write_data[37]));
DFF_X1 \my_reg_reg[38]  (.Q (read_data[38]), .CK (CTS_n_tid1_7), .D (write_data[38]));
DFF_X1 \my_reg_reg[39]  (.Q (read_data[39]), .CK (CTS_n_tid1_7), .D (write_data[39]));
DFF_X1 \my_reg_reg[40]  (.Q (read_data[40]), .CK (CTS_n_tid1_7), .D (write_data[40]));
DFF_X1 \my_reg_reg[41]  (.Q (read_data[41]), .CK (CTS_n_tid1_7), .D (write_data[41]));
DFF_X1 \my_reg_reg[42]  (.Q (read_data[42]), .CK (CTS_n_tid1_7), .D (write_data[42]));
DFF_X1 \my_reg_reg[43]  (.Q (read_data[43]), .CK (CTS_n_tid1_7), .D (write_data[43]));
DFF_X1 \my_reg_reg[44]  (.Q (read_data[44]), .CK (CTS_n_tid1_7), .D (write_data[44]));
DFF_X1 \my_reg_reg[45]  (.Q (read_data[45]), .CK (CTS_n_tid1_7), .D (write_data[45]));
DFF_X1 \my_reg_reg[46]  (.Q (read_data[46]), .CK (CTS_n_tid1_7), .D (write_data[46]));
DFF_X1 \my_reg_reg[47]  (.Q (read_data[47]), .CK (CTS_n_tid1_7), .D (write_data[47]));
DFF_X1 \my_reg_reg[48]  (.Q (read_data[48]), .CK (CTS_n_tid1_7), .D (write_data[48]));
DFF_X1 \my_reg_reg[49]  (.Q (read_data[49]), .CK (CTS_n_tid1_7), .D (write_data[49]));
DFF_X1 \my_reg_reg[50]  (.Q (read_data[50]), .CK (CTS_n_tid1_7), .D (write_data[50]));
DFF_X1 \my_reg_reg[51]  (.Q (read_data[51]), .CK (CTS_n_tid1_7), .D (write_data[51]));
DFF_X1 \my_reg_reg[52]  (.Q (read_data[52]), .CK (CTS_n_tid1_7), .D (write_data[52]));
DFF_X1 \my_reg_reg[53]  (.Q (read_data[53]), .CK (CTS_n_tid1_7), .D (write_data[53]));
DFF_X1 \my_reg_reg[54]  (.Q (read_data[54]), .CK (CTS_n_tid1_7), .D (write_data[54]));
DFF_X1 \my_reg_reg[55]  (.Q (read_data[55]), .CK (CTS_n_tid1_7), .D (write_data[55]));
DFF_X1 \my_reg_reg[56]  (.Q (read_data[56]), .CK (CTS_n_tid1_7), .D (write_data[56]));
DFF_X1 \my_reg_reg[57]  (.Q (read_data[57]), .CK (CTS_n_tid1_7), .D (write_data[57]));
DFF_X1 \my_reg_reg[58]  (.Q (read_data[58]), .CK (CTS_n_tid1_7), .D (write_data[58]));
DFF_X1 \my_reg_reg[59]  (.Q (read_data[59]), .CK (CTS_n_tid1_7), .D (write_data[59]));
DFF_X1 \my_reg_reg[60]  (.Q (read_data[60]), .CK (CTS_n_tid1_7), .D (write_data[60]));
DFF_X1 \my_reg_reg[61]  (.Q (read_data[61]), .CK (CTS_n_tid1_7), .D (write_data[61]));
DFF_X1 \my_reg_reg[62]  (.Q (read_data[62]), .CK (CTS_n_tid1_7), .D (write_data[62]));
CLKBUF_X3 CTS_L3_c_tid1_4 (.Z (CTS_n_tid1_7), .A (n_tid1_34));
DFF_X1 \my_reg_reg[63]  (.Q (read_data[63]), .CK (CTS_n_tid1_7), .D (write_data[63]));
INV_X4 CTS_L2_tid1__c2_tid1__c11 (.ZN (n_tid1_34), .A (clk__CTS_1_PP_1));

endmodule //regFile64

module full_adder (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


XNOR2_X1 i_0_5 (.ZN (n_0_4), .A (i_bit1), .B (i_bit2));
NAND2_X1 i_0_4 (.ZN (n_0_3), .A1 (i_carry), .A2 (n_0_4));
INV_X1 i_0_3 (.ZN (n_0_2), .A (i_carry));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_0 (.ZN (o_sum), .A1 (n_0_0), .A2 (n_0_3));

endmodule //full_adder

module full_adder__0_465 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


XNOR2_X1 i_0_5 (.ZN (n_0_4), .A (i_bit1), .B (i_bit2));
NAND2_X1 i_0_4 (.ZN (n_0_3), .A1 (i_carry), .A2 (n_0_4));
INV_X1 i_0_3 (.ZN (n_0_2), .A (i_carry));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_0 (.ZN (o_sum), .A1 (n_0_0), .A2 (n_0_3));

endmodule //full_adder__0_465

module full_adder__0_461 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_461

module full_adder__0_457 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_457

module full_adder__0_453 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_453

module full_adder__0_449 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_449

module full_adder__0_445 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_445

module full_adder__0_441 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_441

module full_adder__0_437 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_437

module full_adder__0_433 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_433

module full_adder__0_429 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_429

module full_adder__0_425 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_425

module full_adder__0_421 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_421

module full_adder__0_417 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_417

module full_adder__0_413 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_413

module full_adder__0_409 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_409

module full_adder__0_405 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_405

module full_adder__0_401 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_401

module full_adder__0_397 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_397

module full_adder__0_393 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_393

module full_adder__0_389 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_389

module full_adder__0_385 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_385

module full_adder__0_381 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_381

module full_adder__0_377 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_377

module full_adder__0_373 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_373

module full_adder__0_369 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_369

module full_adder__0_365 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_365

module full_adder__0_361 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_361

module full_adder__0_357 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_357

module full_adder__0_353 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_353

module full_adder__0_349 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_349

module full_adder__0_345 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_345

module full_adder__0_341 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_341

module full_adder__0_337 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_337

module full_adder__0_333 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_333

module full_adder__0_329 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_329

module full_adder__0_325 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_325

module full_adder__0_321 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_321

module full_adder__0_317 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_317

module full_adder__0_313 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_313

module full_adder__0_309 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_309

module full_adder__0_305 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_305

module full_adder__0_301 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_301

module full_adder__0_297 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_297

module full_adder__0_293 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_293

module full_adder__0_289 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_289

module full_adder__0_285 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_285

module full_adder__0_281 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_281

module full_adder__0_277 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_277

module full_adder__0_273 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_273

module full_adder__0_269 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_269

module full_adder__0_265 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_265

module full_adder__0_261 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_261

module full_adder__0_257 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_257

module full_adder__0_253 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_253

module full_adder__0_249 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_249

module full_adder__0_245 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_245

module full_adder__0_241 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_241

module full_adder__0_237 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_237

module full_adder__0_233 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_233

module full_adder__0_229 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_229

module full_adder__0_225 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_225

module full_adder__0_221 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;
wire n_0_0;


XOR2_X1 i_0_1 (.Z (o_sum), .A (n_0_0), .B (i_carry));
XOR2_X1 i_0_0 (.Z (n_0_0), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_221

module full_adder__0_217 (i_bit1, i_bit2, i_carry, o_sum, o_carry);

output o_carry;
output o_sum;
input i_bit1;
input i_bit2;
input i_carry;


XOR2_X1 i_0_0 (.Z (o_sum), .A (i_bit1), .B (i_bit2));

endmodule //full_adder__0_217

module carry_lookahead_adder (i_add1, i_add2, o_result, o_carry);

output o_carry;
output [63:0] o_result;
input [63:0] i_add1;
input [63:0] i_add2;
wire n_0_38;
wire n_0_21;
wire n_0_27;
wire n_0_39;
wire n_0_40;
wire n_0_35;
wire n_0_41;
wire n_0_42;
wire w_G;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_155;
wire n_0_157;
wire n_0_47;
wire n_0_168;
wire n_0_48;
wire n_0_201;
wire n_0_202;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_237;
wire n_0_49;
wire n_0_259;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_50;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_51;
wire n_0_384;
wire n_0_385;
wire n_0_386;
wire n_0_387;
wire n_0_388;
wire n_0_181;
wire n_0_389;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_171;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_146;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_111;
wire n_0_19;
wire n_0_101;
wire n_0_20;
wire n_0_22;
wire n_0_96;
wire n_0_23;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_156;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_169;
wire n_0_170;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_214;
wire n_0_215;
wire n_0_217;
wire n_0_218;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_234;
wire n_0_236;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_260;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_296;
wire n_0_297;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_317;
wire n_0_318;
wire n_0_319;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_328;
wire n_0_329;
wire n_0_330;
wire n_0_331;
wire n_0_332;
wire n_0_333;
wire n_0_334;
wire n_0_335;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_339;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_344;
wire n_0_345;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_351;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_355;
wire n_0_356;
wire n_0_357;
wire n_0_358;
wire n_0_359;
wire n_0_360;
wire n_0_361;
wire n_0_362;
wire n_0_363;
wire n_0_365;
wire n_0_366;
wire n_0_367;
wire n_0_368;
wire n_0_369;
wire n_0_370;
wire n_0_372;
wire n_0_373;
wire n_0_374;
wire n_0_375;
wire n_0_376;
wire n_0_377;
wire n_0_378;
wire n_0_379;
wire n_0_380;
wire n_0_381;
wire n_0_382;
wire n_0_383;
wire n_61;
wire n_23;
wire n_60;
wire n_22;
wire n_59;
wire n_21;
wire n_58;
wire n_57;
wire n_56;
wire n_20;
wire n_55;
wire n_19;
wire n_54;
wire n_18;
wire n_53;
wire n_52;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_51;
wire n_10;
wire n_9;
wire n_8;
wire n_50;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire n_42;
wire n_49;
wire n_48;
wire n_47;
wire n_46;


AND2_X1 i_0_422 (.ZN (n_61), .A1 (n_0_379), .A2 (n_0_378));
INV_X1 i_0_421 (.ZN (n_0_383), .A (i_add2[3]));
INV_X1 i_0_420 (.ZN (n_0_382), .A (i_add1[3]));
NAND2_X1 i_0_419 (.ZN (n_0_381), .A1 (i_add2[0]), .A2 (i_add1[0]));
NAND2_X1 i_0_418 (.ZN (n_0_380), .A1 (i_add2[1]), .A2 (i_add1[1]));
NAND2_X1 i_0_417 (.ZN (n_0_379), .A1 (n_0_381), .A2 (n_0_380));
OR2_X1 i_0_416 (.ZN (n_0_378), .A1 (i_add2[1]), .A2 (i_add1[1]));
AOI22_X1 i_0_415 (.ZN (n_0_377), .A1 (n_0_379), .A2 (n_0_378), .B1 (i_add2[2]), .B2 (i_add1[2]));
NOR2_X1 i_0_414 (.ZN (n_0_376), .A1 (i_add2[2]), .A2 (i_add1[2]));
OAI22_X1 i_0_413 (.ZN (n_0_375), .A1 (n_0_383), .A2 (n_0_382), .B1 (n_0_377), .B2 (n_0_376));
NAND2_X1 i_0_412 (.ZN (n_0_374), .A1 (n_0_383), .A2 (n_0_382));
AND2_X1 i_0_411 (.ZN (n_60), .A1 (n_0_375), .A2 (n_0_374));
AND2_X1 i_0_410 (.ZN (n_0_373), .A1 (i_add2[4]), .A2 (i_add1[4]));
AND2_X1 i_0_409 (.ZN (n_59), .A1 (n_0_222), .A2 (n_0_208));
AND2_X1 i_0_408 (.ZN (n_58), .A1 (n_0_366), .A2 (n_0_210));
INV_X1 i_0_407 (.ZN (n_0_372), .A (n_0_214));
AND2_X1 i_0_405 (.ZN (n_0_370), .A1 (i_add1[8]), .A2 (i_add2[8]));
NAND2_X1 i_0_404 (.ZN (n_0_369), .A1 (i_add1[7]), .A2 (i_add2[7]));
AND2_X1 i_0_403 (.ZN (n_0_368), .A1 (i_add1[6]), .A2 (i_add2[6]));
AOI21_X1 i_0_402 (.ZN (n_0_367), .A (n_0_368), .B1 (n_0_222), .B2 (n_0_208));
OAI21_X1 i_0_401 (.ZN (n_0_366), .A (n_0_369), .B1 (n_0_372), .B2 (n_0_367));
AOI21_X1 i_0_400 (.ZN (n_0_365), .A (n_0_370), .B1 (n_0_210), .B2 (n_0_366));
NOR2_X1 i_0_399 (.ZN (n_57), .A1 (n_0_212), .A2 (n_0_365));
AND2_X1 i_0_398 (.ZN (n_56), .A1 (n_0_357), .A2 (n_0_356));
AOI21_X1 i_0_396 (.ZN (n_0_363), .A (n_0_347), .B1 (n_0_356), .B2 (n_0_357));
OAI21_X1 i_0_395 (.ZN (n_0_362), .A (n_0_205), .B1 (n_0_340), .B2 (n_0_363));
AND2_X1 i_0_394 (.ZN (n_55), .A1 (n_0_355), .A2 (n_0_362));
INV_X1 i_0_393 (.ZN (n_0_361), .A (i_add1[11]));
INV_X1 i_0_392 (.ZN (n_0_360), .A (i_add2[11]));
INV_X1 i_0_391 (.ZN (n_0_359), .A (n_0_221));
INV_X1 i_0_390 (.ZN (n_0_358), .A (n_0_341));
NAND2_X1 i_0_389 (.ZN (n_0_357), .A1 (n_0_343), .A2 (n_0_204));
OR2_X1 i_0_388 (.ZN (n_0_356), .A1 (i_add1[9]), .A2 (i_add2[9]));
NAND2_X1 i_0_387 (.ZN (n_0_355), .A1 (n_0_361), .A2 (n_0_360));
AOI21_X1 i_0_386 (.ZN (n_0_354), .A (n_0_347), .B1 (n_0_357), .B2 (n_0_356));
OAI21_X1 i_0_385 (.ZN (n_0_353), .A (n_0_205), .B1 (n_0_340), .B2 (n_0_354));
AOI21_X1 i_0_384 (.ZN (n_0_352), .A (n_0_359), .B1 (n_0_355), .B2 (n_0_353));
OAI21_X1 i_0_383 (.ZN (n_0_351), .A (n_0_336), .B1 (n_0_358), .B2 (n_0_352));
AND2_X1 i_0_382 (.ZN (n_54), .A1 (n_0_215), .A2 (n_0_351));
AOI21_X1 i_0_380 (.ZN (n_0_349), .A (n_0_344), .B1 (n_0_334), .B2 (n_0_215));
OAI21_X1 i_0_379 (.ZN (n_0_348), .A (n_0_187), .B1 (n_0_333), .B2 (n_0_349));
AND2_X1 i_0_378 (.ZN (n_53), .A1 (n_0_346), .A2 (n_0_348));
INV_X1 i_0_377 (.ZN (n_0_347), .A (n_0_206));
INV_X1 i_0_376 (.ZN (n_0_346), .A (n_0_188));
NAND2_X1 i_0_375 (.ZN (n_0_345), .A1 (i_add2[14]), .A2 (i_add1[14]));
INV_X1 i_0_374 (.ZN (n_0_344), .A (n_0_345));
AOI21_X1 i_0_373 (.ZN (n_0_343), .A (n_0_198), .B1 (n_0_222), .B2 (n_0_207));
INV_X1 i_0_372 (.ZN (n_0_342), .A (n_0_343));
OR2_X1 i_0_371 (.ZN (n_0_341), .A1 (i_add2[12]), .A2 (i_add1[12]));
NOR2_X1 i_0_370 (.ZN (n_0_340), .A1 (i_add2[10]), .A2 (i_add1[10]));
NOR3_X1 i_0_369 (.ZN (n_0_339), .A1 (i_add2[9]), .A2 (n_0_347), .A3 (i_add1[9]));
OAI211_X1 i_0_368 (.ZN (n_0_338), .A (n_0_205), .B (n_0_221), .C1 (n_0_340), .C2 (n_0_339));
INV_X1 i_0_367 (.ZN (n_0_337), .A (n_0_338));
NAND2_X1 i_0_366 (.ZN (n_0_336), .A1 (i_add2[13]), .A2 (i_add1[13]));
OAI211_X1 i_0_365 (.ZN (n_0_335), .A (n_0_220), .B (n_0_341), .C1 (n_0_203), .C2 (n_0_342));
OAI21_X1 i_0_364 (.ZN (n_0_334), .A (n_0_336), .B1 (n_0_337), .B2 (n_0_335));
NOR2_X1 i_0_363 (.ZN (n_0_333), .A1 (i_add2[14]), .A2 (i_add1[14]));
INV_X1 i_0_362 (.ZN (n_0_332), .A (n_0_333));
NAND3_X1 i_0_361 (.ZN (n_0_331), .A1 (n_0_215), .A2 (n_0_332), .A3 (n_0_334));
NAND2_X1 i_0_360 (.ZN (n_0_330), .A1 (n_0_187), .A2 (n_0_331));
OAI21_X1 i_0_359 (.ZN (n_0_329), .A (n_0_346), .B1 (n_0_344), .B2 (n_0_330));
AOI21_X1 i_0_358 (.ZN (n_52), .A (n_0_257), .B1 (n_0_179), .B2 (n_0_329));
AOI21_X1 i_0_357 (.ZN (n_0_328), .A (n_0_228), .B1 (n_0_245), .B2 (n_0_158));
INV_X1 i_0_356 (.ZN (n_0_327), .A (n_0_328));
AOI21_X1 i_0_355 (.ZN (n_51), .A (n_0_105), .B1 (n_0_159), .B2 (n_0_327));
INV_X1 i_0_354 (.ZN (n_0_326), .A (n_51));
NOR2_X1 i_0_353 (.ZN (n_0_325), .A1 (n_0_240), .A2 (n_0_129));
NOR2_X1 i_0_352 (.ZN (n_50), .A1 (n_0_88), .A2 (n_0_325));
OR2_X1 i_0_351 (.ZN (n_49), .A1 (n_0_282), .A2 (n_0_279));
NOR3_X1 i_0_350 (.ZN (n_0_324), .A1 (n_0_279), .A2 (n_0_277), .A3 (n_0_282));
NOR2_X1 i_0_349 (.ZN (n_0_323), .A1 (n_0_273), .A2 (n_0_324));
NOR2_X1 i_0_348 (.ZN (n_0_322), .A1 (n_0_278), .A2 (n_0_323));
NOR2_X1 i_0_347 (.ZN (n_48), .A1 (n_0_274), .A2 (n_0_322));
AOI21_X1 i_0_346 (.ZN (n_47), .A (n_0_320), .B1 (n_0_321), .B2 (n_0_307));
INV_X1 i_0_345 (.ZN (n_0_321), .A (n_0_319));
INV_X1 i_0_344 (.ZN (n_0_320), .A (n_0_270));
AOI221_X1 i_0_343 (.ZN (n_0_319), .A (n_0_271), .B1 (n_0_315), .B2 (n_0_316), .C1 (n_0_318), .C2 (n_0_316));
NOR3_X1 i_0_342 (.ZN (n_0_318), .A1 (n_0_317), .A2 (n_0_58), .A3 (n_0_303));
AND3_X1 i_0_341 (.ZN (n_0_317), .A1 (n_0_99), .A2 (n_0_69), .A3 (n_0_124));
NOR2_X1 i_0_340 (.ZN (n_0_316), .A1 (n_0_279), .A2 (n_0_275));
OR2_X1 i_0_339 (.ZN (n_0_315), .A1 (n_0_283), .A2 (n_0_287));
INV_X1 i_0_338 (.ZN (n_0_314), .A (i_add2[58]));
INV_X1 i_0_337 (.ZN (n_0_313), .A (i_add2[57]));
INV_X1 i_0_336 (.ZN (n_0_312), .A (i_add2[55]));
INV_X1 i_0_335 (.ZN (n_0_311), .A (i_add1[58]));
INV_X1 i_0_334 (.ZN (n_0_310), .A (i_add1[57]));
INV_X1 i_0_333 (.ZN (n_0_309), .A (i_add1[55]));
INV_X1 i_0_332 (.ZN (n_0_308), .A (n_0_53));
NAND2_X1 i_0_331 (.ZN (n_0_307), .A1 (i_add2[61]), .A2 (i_add1[61]));
INV_X1 i_0_330 (.ZN (n_0_306), .A (n_0_307));
NAND2_X1 i_0_329 (.ZN (n_0_305), .A1 (i_add2[53]), .A2 (i_add1[53]));
AOI21_X1 i_0_328 (.ZN (n_0_304), .A (n_0_308), .B1 (i_add2[54]), .B2 (i_add1[54]));
NAND3_X1 i_0_327 (.ZN (n_0_303), .A1 (n_0_56), .A2 (n_0_305), .A3 (n_0_304));
INV_X1 i_0_326 (.ZN (n_0_302), .A (n_0_303));
NAND3_X1 i_0_325 (.ZN (n_0_297), .A1 (n_0_68), .A2 (n_0_302), .A3 (n_0_59));
INV_X1 i_0_324 (.ZN (n_0_296), .A (n_0_297));
OR2_X1 i_0_323 (.ZN (n_0_292), .A1 (i_add2[54]), .A2 (i_add1[54]));
NAND2_X1 i_0_322 (.ZN (n_0_291), .A1 (n_0_312), .A2 (n_0_309));
NOR2_X1 i_0_321 (.ZN (n_0_290), .A1 (i_add2[56]), .A2 (i_add1[56]));
AOI21_X1 i_0_320 (.ZN (n_0_289), .A (n_0_290), .B1 (n_0_313), .B2 (n_0_310));
INV_X1 i_0_319 (.ZN (n_0_288), .A (n_0_289));
NAND3_X1 i_0_318 (.ZN (n_0_287), .A1 (n_0_292), .A2 (n_0_291), .A3 (n_0_289));
OR2_X1 i_0_317 (.ZN (n_0_286), .A1 (i_add2[53]), .A2 (i_add1[53]));
NOR3_X1 i_0_316 (.ZN (n_0_285), .A1 (i_add2[51]), .A2 (n_0_308), .A3 (i_add1[51]));
OAI21_X1 i_0_315 (.ZN (n_0_284), .A (n_0_305), .B1 (n_0_226), .B2 (n_0_285));
AOI22_X1 i_0_314 (.ZN (n_0_283), .A1 (i_add2[54]), .A2 (i_add1[54]), .B1 (n_0_286), .B2 (n_0_284));
NOR3_X1 i_0_313 (.ZN (n_0_282), .A1 (n_0_287), .A2 (n_0_283), .A3 (n_0_296));
NOR2_X1 i_0_312 (.ZN (n_0_281), .A1 (n_0_312), .A2 (n_0_309));
AOI21_X1 i_0_311 (.ZN (n_0_280), .A (n_0_281), .B1 (i_add2[56]), .B2 (i_add1[56]));
OAI22_X1 i_0_310 (.ZN (n_0_279), .A1 (n_0_313), .A2 (n_0_310), .B1 (n_0_288), .B2 (n_0_280));
AND2_X1 i_0_309 (.ZN (n_0_278), .A1 (i_add2[59]), .A2 (i_add1[59]));
NOR2_X1 i_0_308 (.ZN (n_0_277), .A1 (n_0_314), .A2 (n_0_311));
AOI21_X1 i_0_307 (.ZN (n_0_276), .A (n_0_278), .B1 (i_add2[60]), .B2 (i_add1[60]));
OAI21_X1 i_0_306 (.ZN (n_0_275), .A (n_0_276), .B1 (n_0_314), .B2 (n_0_311));
NOR2_X1 i_0_305 (.ZN (n_0_274), .A1 (i_add2[59]), .A2 (i_add1[59]));
NOR2_X1 i_0_304 (.ZN (n_0_273), .A1 (i_add2[58]), .A2 (i_add1[58]));
OAI21_X1 i_0_303 (.ZN (n_0_272), .A (n_0_276), .B1 (n_0_274), .B2 (n_0_273));
OAI21_X1 i_0_302 (.ZN (n_0_271), .A (n_0_272), .B1 (i_add2[60]), .B2 (i_add1[60]));
OR2_X1 i_0_301 (.ZN (n_0_270), .A1 (i_add2[61]), .A2 (i_add1[61]));
NAND2_X1 i_0_300 (.ZN (n_0_269), .A1 (i_add2[62]), .A2 (i_add1[62]));
NOR3_X1 i_0_299 (.ZN (n_0_268), .A1 (n_0_282), .A2 (n_0_279), .A3 (n_0_275));
NOR2_X1 i_0_298 (.ZN (n_0_267), .A1 (n_0_271), .A2 (n_0_268));
OAI221_X1 i_0_297 (.ZN (n_0_266), .A (n_0_270), .B1 (i_add2[62]), .B2 (i_add1[62])
    , .C1 (n_0_306), .C2 (n_0_267));
NAND2_X1 i_0_296 (.ZN (n_46), .A1 (n_0_269), .A2 (n_0_266));
INV_X1 i_0_295 (.ZN (n_0_265), .A (n_0_179));
NOR2_X1 i_0_294 (.ZN (n_0_260), .A1 (i_add2[18]), .A2 (i_add1[18]));
INV_X1 i_0_293 (.ZN (n_0_258), .A (n_0_260));
NOR2_X1 i_0_292 (.ZN (n_0_257), .A1 (i_add2[16]), .A2 (i_add1[16]));
INV_X1 i_0_291 (.ZN (n_0_256), .A (n_0_257));
OR2_X1 i_0_290 (.ZN (n_0_255), .A1 (i_add2[17]), .A2 (i_add1[17]));
NOR3_X1 i_0_289 (.ZN (n_0_254), .A1 (n_0_265), .A2 (n_0_195), .A3 (n_0_184));
OAI21_X1 i_0_288 (.ZN (n_0_253), .A (n_0_177), .B1 (n_0_257), .B2 (n_0_254));
NAND2_X1 i_0_287 (.ZN (n_0_252), .A1 (n_0_255), .A2 (n_0_253));
AOI21_X1 i_0_286 (.ZN (n_0_251), .A (n_0_260), .B1 (n_0_175), .B2 (n_0_252));
INV_X1 i_0_285 (.ZN (n_0_250), .A (n_0_89));
INV_X1 i_0_283 (.ZN (n_0_248), .A (n_0_149));
NOR2_X1 i_0_282 (.ZN (n_0_247), .A1 (n_0_195), .A2 (n_0_165));
NOR2_X1 i_0_281 (.ZN (n_0_246), .A1 (n_0_134), .A2 (n_0_247));
AOI21_X1 i_0_280 (.ZN (n_0_245), .A (n_0_160), .B1 (n_0_117), .B2 (n_0_246));
NAND2_X1 i_0_279 (.ZN (n_0_244), .A1 (n_0_150), .A2 (n_0_245));
NAND3_X1 i_0_278 (.ZN (n_0_243), .A1 (n_0_102), .A2 (n_0_244), .A3 (n_0_108));
NAND2_X1 i_0_277 (.ZN (n_0_242), .A1 (n_0_164), .A2 (n_0_243));
OAI22_X1 i_0_276 (.ZN (n_0_241), .A1 (i_add2[37]), .A2 (i_add1[37]), .B1 (n_0_248), .B2 (n_0_242));
AOI21_X1 i_0_275 (.ZN (n_0_240), .A (n_0_250), .B1 (n_0_148), .B2 (n_0_241));
INV_X1 i_0_274 (.ZN (n_0_239), .A (i_add2[43]));
INV_X1 i_0_273 (.ZN (n_0_236), .A (i_add1[43]));
INV_X1 i_0_272 (.ZN (n_0_234), .A (n_0_42));
INV_X1 i_0_271 (.ZN (n_0_229), .A (n_0_50));
INV_X1 i_0_270 (.ZN (n_0_228), .A (n_0_39));
INV_X1 i_0_269 (.ZN (n_0_227), .A (n_0_38));
NOR2_X1 i_0_268 (.ZN (n_0_226), .A1 (i_add2[52]), .A2 (i_add1[52]));
AOI21_X1 i_0_267 (.ZN (n_0_225), .A (n_0_373), .B1 (n_0_375), .B2 (n_0_374));
NAND2_X1 i_0_266 (.ZN (n_0_224), .A1 (i_add2[5]), .A2 (i_add1[5]));
OAI21_X1 i_0_265 (.ZN (n_0_222), .A (n_0_224), .B1 (n_0_234), .B2 (n_0_225));
NAND2_X1 i_0_264 (.ZN (n_0_221), .A1 (i_add2[12]), .A2 (i_add1[12]));
NAND3_X1 i_0_263 (.ZN (n_0_220), .A1 (n_0_360), .A2 (n_0_221), .A3 (n_0_361));
INV_X1 i_0_262 (.ZN (n_0_218), .A (n_0_220));
NOR2_X1 i_0_261 (.ZN (n_0_217), .A1 (i_add2[13]), .A2 (i_add1[13]));
INV_X1 i_0_260 (.ZN (n_0_215), .A (n_0_217));
OR2_X1 i_0_259 (.ZN (n_0_214), .A1 (i_add2[6]), .A2 (i_add1[6]));
NOR2_X1 i_0_258 (.ZN (n_0_212), .A1 (i_add2[8]), .A2 (i_add1[8]));
INV_X1 i_0_257 (.ZN (n_0_211), .A (n_0_212));
OR2_X1 i_0_256 (.ZN (n_0_210), .A1 (i_add2[7]), .A2 (i_add1[7]));
OR2_X1 i_0_255 (.ZN (n_0_208), .A1 (i_add2[5]), .A2 (i_add1[5]));
AND4_X1 i_0_254 (.ZN (n_0_207), .A1 (n_0_214), .A2 (n_0_211), .A3 (n_0_210), .A4 (n_0_208));
NAND2_X1 i_0_253 (.ZN (n_0_206), .A1 (i_add2[10]), .A2 (i_add1[10]));
NAND2_X1 i_0_252 (.ZN (n_0_205), .A1 (i_add2[11]), .A2 (i_add1[11]));
NAND2_X1 i_0_251 (.ZN (n_0_204), .A1 (i_add2[9]), .A2 (i_add1[9]));
NAND4_X1 i_0_250 (.ZN (n_0_203), .A1 (n_0_221), .A2 (n_0_206), .A3 (n_0_205), .A4 (n_0_204));
NOR2_X1 i_0_249 (.ZN (n_0_200), .A1 (n_0_370), .A2 (n_0_44));
NAND3_X1 i_0_248 (.ZN (n_0_199), .A1 (n_0_214), .A2 (n_0_210), .A3 (n_0_368));
AOI21_X1 i_0_247 (.ZN (n_0_198), .A (n_0_212), .B1 (n_0_200), .B2 (n_0_199));
AOI211_X1 i_0_246 (.ZN (n_0_197), .A (n_0_203), .B (n_0_198), .C1 (n_0_222), .C2 (n_0_207));
NAND4_X1 i_0_245 (.ZN (n_0_196), .A1 (n_0_338), .A2 (n_0_346), .A3 (n_0_332), .A4 (n_0_341));
NOR4_X1 i_0_244 (.ZN (n_0_195), .A1 (n_0_217), .A2 (n_0_196), .A3 (n_0_218), .A4 (n_0_197));
OR2_X1 i_0_243 (.ZN (n_0_194), .A1 (i_add2[21]), .A2 (i_add1[21]));
NOR2_X1 i_0_242 (.ZN (n_0_193), .A1 (i_add2[22]), .A2 (i_add1[22]));
INV_X1 i_0_241 (.ZN (n_0_192), .A (n_0_193));
AND2_X1 i_0_240 (.ZN (n_0_190), .A1 (n_0_48), .A2 (n_0_194));
AOI22_X1 i_0_239 (.ZN (n_0_189), .A1 (i_add2[22]), .A2 (i_add1[22]), .B1 (n_0_192), .B2 (n_0_190));
NOR2_X1 i_0_238 (.ZN (n_0_188), .A1 (i_add2[15]), .A2 (i_add1[15]));
NAND2_X1 i_0_237 (.ZN (n_0_187), .A1 (i_add2[15]), .A2 (i_add1[15]));
OAI21_X1 i_0_236 (.ZN (n_0_185), .A (n_0_332), .B1 (n_0_344), .B2 (n_0_45));
OAI21_X1 i_0_235 (.ZN (n_0_184), .A (n_0_187), .B1 (n_0_188), .B2 (n_0_185));
AND2_X1 i_0_234 (.ZN (n_0_183), .A1 (i_add2[23]), .A2 (i_add1[23]));
AND2_X1 i_0_233 (.ZN (n_0_182), .A1 (i_add2[25]), .A2 (i_add1[25]));
NAND2_X1 i_0_232 (.ZN (n_0_180), .A1 (i_add2[24]), .A2 (i_add1[24]));
NAND2_X1 i_0_231 (.ZN (n_0_179), .A1 (i_add2[16]), .A2 (i_add1[16]));
NAND2_X1 i_0_230 (.ZN (n_0_178), .A1 (i_add2[19]), .A2 (i_add1[19]));
NAND2_X1 i_0_229 (.ZN (n_0_177), .A1 (i_add2[17]), .A2 (i_add1[17]));
NAND2_X1 i_0_228 (.ZN (n_0_175), .A1 (i_add2[18]), .A2 (i_add1[18]));
NAND4_X1 i_0_227 (.ZN (n_0_174), .A1 (n_0_179), .A2 (n_0_178), .A3 (n_0_177), .A4 (n_0_175));
AND2_X1 i_0_226 (.ZN (n_0_173), .A1 (i_add2[26]), .A2 (i_add1[26]));
NOR2_X1 i_0_225 (.ZN (n_0_172), .A1 (n_0_183), .A2 (n_0_173));
AOI21_X1 i_0_224 (.ZN (n_0_170), .A (n_0_182), .B1 (i_add2[24]), .B2 (i_add1[24]));
NAND3_X1 i_0_223 (.ZN (n_0_169), .A1 (n_0_172), .A2 (n_0_170), .A3 (n_0_189));
OR3_X1 i_0_222 (.ZN (n_0_165), .A1 (n_0_184), .A2 (n_0_174), .A3 (n_0_169));
OAI21_X1 i_0_221 (.ZN (n_0_164), .A (n_0_229), .B1 (i_add2[36]), .B2 (i_add1[36]));
NOR2_X1 i_0_220 (.ZN (n_0_163), .A1 (i_add2[29]), .A2 (i_add1[29]));
INV_X1 i_0_219 (.ZN (n_0_162), .A (n_0_163));
AOI21_X1 i_0_218 (.ZN (n_0_160), .A (n_0_163), .B1 (n_0_49), .B2 (n_0_40));
NAND2_X1 i_0_217 (.ZN (n_0_159), .A1 (i_add2[31]), .A2 (i_add1[31]));
NAND2_X1 i_0_216 (.ZN (n_0_158), .A1 (i_add2[30]), .A2 (i_add1[30]));
NAND2_X1 i_0_215 (.ZN (n_0_156), .A1 (i_add2[32]), .A2 (i_add1[32]));
AND2_X1 i_0_214 (.ZN (n_0_154), .A1 (n_0_159), .A2 (n_0_156));
NAND2_X1 i_0_213 (.ZN (n_0_153), .A1 (i_add2[33]), .A2 (i_add1[33]));
NAND3_X1 i_0_212 (.ZN (n_0_152), .A1 (n_0_158), .A2 (n_0_153), .A3 (n_0_154));
INV_X1 i_0_211 (.ZN (n_0_150), .A (n_0_152));
NAND2_X1 i_0_210 (.ZN (n_0_149), .A1 (i_add2[37]), .A2 (i_add1[37]));
NAND2_X1 i_0_209 (.ZN (n_0_148), .A1 (i_add2[38]), .A2 (i_add1[38]));
AOI21_X1 i_0_208 (.ZN (n_0_147), .A (n_0_46), .B1 (n_0_47), .B2 (n_0_258));
NOR2_X1 i_0_207 (.ZN (n_0_145), .A1 (i_add2[20]), .A2 (i_add1[20]));
INV_X1 i_0_206 (.ZN (n_0_144), .A (n_0_145));
OR2_X1 i_0_205 (.ZN (n_0_143), .A1 (i_add2[19]), .A2 (i_add1[19]));
NAND2_X1 i_0_204 (.ZN (n_0_142), .A1 (n_0_194), .A2 (n_0_143));
INV_X1 i_0_203 (.ZN (n_0_140), .A (n_0_142));
NOR2_X1 i_0_202 (.ZN (n_0_139), .A1 (i_add2[25]), .A2 (i_add1[25]));
OR2_X1 i_0_201 (.ZN (n_0_138), .A1 (i_add2[24]), .A2 (i_add1[24]));
NOR4_X1 i_0_200 (.ZN (n_0_137), .A1 (n_0_147), .A2 (n_0_145), .A3 (n_0_142), .A4 (n_0_193));
OAI21_X1 i_0_199 (.ZN (n_0_136), .A (n_0_138), .B1 (i_add2[23]), .B2 (i_add1[23]));
AOI21_X1 i_0_198 (.ZN (n_0_135), .A (n_0_139), .B1 (n_0_170), .B2 (n_0_136));
OAI22_X1 i_0_197 (.ZN (n_0_134), .A1 (n_0_169), .A2 (n_0_137), .B1 (n_0_173), .B2 (n_0_135));
NOR2_X1 i_0_196 (.ZN (n_0_133), .A1 (n_0_195), .A2 (n_0_165));
NOR2_X1 i_0_195 (.ZN (n_0_132), .A1 (n_0_160), .A2 (n_0_152));
INV_X1 i_0_194 (.ZN (n_0_130), .A (n_0_132));
AND2_X1 i_0_193 (.ZN (n_0_129), .A1 (i_add2[39]), .A2 (i_add1[39]));
AOI21_X1 i_0_192 (.ZN (n_0_128), .A (n_0_129), .B1 (i_add2[38]), .B2 (i_add1[38]));
NAND2_X1 i_0_191 (.ZN (n_0_127), .A1 (i_add2[40]), .A2 (i_add1[40]));
AND4_X1 i_0_190 (.ZN (n_0_125), .A1 (n_0_149), .A2 (n_0_127), .A3 (n_0_164), .A4 (n_0_128));
OAI211_X1 i_0_189 (.ZN (n_0_124), .A (n_0_132), .B (n_0_125), .C1 (n_0_134), .C2 (n_0_133));
OR2_X1 i_0_187 (.ZN (n_0_123), .A1 (i_add2[26]), .A2 (i_add1[26]));
OR2_X1 i_0_186 (.ZN (n_0_122), .A1 (i_add2[28]), .A2 (i_add1[28]));
NOR2_X1 i_0_185 (.ZN (n_0_120), .A1 (i_add2[27]), .A2 (i_add1[27]));
INV_X1 i_0_184 (.ZN (n_0_119), .A (n_0_120));
NAND4_X1 i_0_183 (.ZN (n_0_118), .A1 (n_0_123), .A2 (n_0_122), .A3 (n_0_119), .A4 (n_0_162));
INV_X1 i_0_182 (.ZN (n_0_117), .A (n_0_118));
OR2_X1 i_0_181 (.ZN (n_0_115), .A1 (i_add2[34]), .A2 (i_add1[34]));
NOR2_X1 i_0_180 (.ZN (n_0_114), .A1 (i_add2[35]), .A2 (i_add1[35]));
INV_X1 i_0_179 (.ZN (n_0_113), .A (n_0_114));
NOR2_X1 i_0_178 (.ZN (n_0_112), .A1 (i_add2[33]), .A2 (i_add1[33]));
INV_X1 i_0_177 (.ZN (n_0_110), .A (n_0_112));
OAI21_X1 i_0_175 (.ZN (n_0_109), .A (n_0_115), .B1 (i_add2[36]), .B2 (i_add1[36]));
NOR3_X1 i_0_174 (.ZN (n_0_108), .A1 (n_0_114), .A2 (n_0_109), .A3 (n_0_112));
OR2_X1 i_0_173 (.ZN (n_0_107), .A1 (i_add2[32]), .A2 (i_add1[32]));
NOR2_X1 i_0_172 (.ZN (n_0_105), .A1 (i_add2[31]), .A2 (i_add1[31]));
OAI21_X1 i_0_171 (.ZN (n_0_104), .A (n_0_154), .B1 (n_0_228), .B2 (n_0_105));
NAND2_X1 i_0_170 (.ZN (n_0_103), .A1 (n_0_107), .A2 (n_0_104));
NAND2_X1 i_0_169 (.ZN (n_0_102), .A1 (n_0_153), .A2 (n_0_103));
OAI211_X1 i_0_168 (.ZN (n_0_100), .A (n_0_108), .B (n_0_102), .C1 (n_0_130), .C2 (n_0_117));
NAND2_X1 i_0_167 (.ZN (n_0_99), .A1 (n_0_125), .A2 (n_0_100));
OR2_X1 i_0_165 (.ZN (n_0_98), .A1 (i_add2[46]), .A2 (i_add1[46]));
NOR2_X1 i_0_164 (.ZN (n_0_97), .A1 (i_add2[45]), .A2 (i_add1[45]));
NAND2_X1 i_0_163 (.ZN (n_0_95), .A1 (i_add2[46]), .A2 (i_add1[46]));
NAND2_X1 i_0_162 (.ZN (n_0_94), .A1 (i_add2[47]), .A2 (i_add1[47]));
NOR2_X1 i_0_161 (.ZN (n_0_93), .A1 (i_add2[48]), .A2 (i_add1[48]));
NOR2_X1 i_0_160 (.ZN (n_0_92), .A1 (i_add2[49]), .A2 (i_add1[49]));
INV_X1 i_0_158 (.ZN (n_0_91), .A (n_0_92));
OR2_X1 i_0_157 (.ZN (n_0_90), .A1 (i_add2[47]), .A2 (i_add1[47]));
OR2_X1 i_0_156 (.ZN (n_0_89), .A1 (i_add2[38]), .A2 (i_add1[38]));
NOR2_X1 i_0_155 (.ZN (n_0_88), .A1 (i_add2[39]), .A2 (i_add1[39]));
OAI21_X1 i_0_154 (.ZN (n_0_87), .A (n_0_89), .B1 (i_add2[37]), .B2 (i_add1[37]));
AOI21_X1 i_0_153 (.ZN (n_0_86), .A (n_0_88), .B1 (n_0_128), .B2 (n_0_87));
AOI21_X1 i_0_152 (.ZN (n_0_85), .A (n_0_86), .B1 (i_add2[40]), .B2 (i_add1[40]));
INV_X1 i_0_151 (.ZN (n_0_84), .A (n_0_85));
OR2_X1 i_0_150 (.ZN (n_0_83), .A1 (i_add2[40]), .A2 (i_add1[40]));
OR2_X1 i_0_149 (.ZN (n_0_82), .A1 (i_add2[42]), .A2 (i_add1[42]));
NOR2_X1 i_0_148 (.ZN (n_0_81), .A1 (i_add2[41]), .A2 (i_add1[41]));
INV_X1 i_0_147 (.ZN (n_0_80), .A (n_0_81));
NOR2_X1 i_0_146 (.ZN (n_0_79), .A1 (i_add2[43]), .A2 (i_add1[43]));
INV_X1 i_0_145 (.ZN (n_0_78), .A (n_0_79));
NAND4_X1 i_0_144 (.ZN (n_0_77), .A1 (n_0_83), .A2 (n_0_82), .A3 (n_0_80), .A4 (n_0_78));
AND2_X1 i_0_143 (.ZN (n_0_76), .A1 (i_add2[45]), .A2 (i_add1[45]));
AOI21_X1 i_0_142 (.ZN (n_0_75), .A (n_0_76), .B1 (i_add2[46]), .B2 (i_add1[46]));
OAI21_X1 i_0_141 (.ZN (n_0_74), .A (n_0_75), .B1 (n_0_227), .B2 (n_0_97));
NAND2_X1 i_0_140 (.ZN (n_0_73), .A1 (n_0_98), .A2 (n_0_74));
NOR2_X1 i_0_139 (.ZN (n_0_72), .A1 (i_add2[50]), .A2 (i_add1[50]));
AOI211_X1 i_0_138 (.ZN (n_0_71), .A (n_0_93), .B (n_0_72), .C1 (n_0_94), .C2 (n_0_73));
NAND3_X1 i_0_137 (.ZN (n_0_70), .A1 (n_0_91), .A2 (n_0_90), .A3 (n_0_71));
NOR3_X1 i_0_136 (.ZN (n_0_69), .A1 (n_0_85), .A2 (n_0_70), .A3 (n_0_77));
NAND3_X1 i_0_135 (.ZN (n_0_68), .A1 (n_0_124), .A2 (n_0_99), .A3 (n_0_69));
NAND2_X1 i_0_134 (.ZN (n_0_67), .A1 (n_0_51), .A2 (n_0_82));
OAI22_X1 i_0_133 (.ZN (n_0_66), .A1 (n_0_239), .A2 (n_0_236), .B1 (n_0_79), .B2 (n_0_67));
NAND2_X1 i_0_132 (.ZN (n_0_65), .A1 (i_add2[44]), .A2 (i_add1[44]));
NAND2_X1 i_0_131 (.ZN (n_0_64), .A1 (i_add2[49]), .A2 (i_add1[49]));
NAND2_X1 i_0_130 (.ZN (n_0_63), .A1 (i_add2[48]), .A2 (i_add1[48]));
AOI221_X1 i_0_129 (.ZN (n_0_62), .A (n_0_66), .B1 (i_add2[47]), .B2 (i_add1[47]), .C1 (i_add2[44]), .C2 (i_add1[44]));
AOI21_X1 i_0_128 (.ZN (n_0_61), .A (n_0_70), .B1 (n_0_75), .B2 (n_0_62));
AOI211_X1 i_0_127 (.ZN (n_0_60), .A (n_0_92), .B (n_0_72), .C1 (n_0_64), .C2 (n_0_63));
AOI211_X1 i_0_126 (.ZN (n_0_59), .A (n_0_61), .B (n_0_60), .C1 (i_add2[50]), .C2 (i_add1[50]));
INV_X1 i_0_125 (.ZN (n_0_58), .A (n_0_59));
NAND2_X1 i_0_124 (.ZN (n_0_57), .A1 (n_0_68), .A2 (n_0_59));
NAND2_X1 i_0_123 (.ZN (n_0_56), .A1 (i_add2[51]), .A2 (i_add1[51]));
INV_X1 i_0_122 (.ZN (n_0_55), .A (n_0_56));
OAI22_X1 i_0_121 (.ZN (n_0_54), .A1 (i_add2[51]), .A2 (i_add1[51]), .B1 (n_0_57), .B2 (n_0_55));
NAND2_X1 i_0_120 (.ZN (n_0_53), .A1 (i_add2[52]), .A2 (i_add1[52]));
AOI21_X1 i_0_119 (.ZN (n_0_52), .A (n_0_226), .B1 (n_0_54), .B2 (n_0_53));
AOI21_X1 i_0_93 (.ZN (n_42), .A (n_0_290), .B1 (n_0_23), .B2 (n_0_280));
NAND4_X1 i_0_92 (.ZN (n_0_23), .A1 (n_0_297), .A2 (n_0_292), .A3 (n_0_291), .A4 (n_0_20));
OAI21_X1 i_0_90 (.ZN (n_0_96), .A (n_0_291), .B1 (n_0_22), .B2 (n_0_281));
AND3_X1 i_0_88 (.ZN (n_0_22), .A1 (n_0_297), .A2 (n_0_292), .A3 (n_0_20));
INV_X1 i_0_87 (.ZN (n_0_20), .A (n_0_283));
OAI21_X1 i_0_86 (.ZN (n_0_101), .A (n_0_286), .B1 (n_0_52), .B2 (n_0_19));
INV_X1 i_0_85 (.ZN (n_0_19), .A (n_0_305));
OAI21_X1 i_0_84 (.ZN (n_0_111), .A (n_0_91), .B1 (n_0_17), .B2 (n_0_18));
INV_X1 i_0_83 (.ZN (n_0_18), .A (n_0_64));
AOI21_X1 i_0_82 (.ZN (n_0_17), .A (n_0_93), .B1 (n_0_16), .B2 (n_0_63));
OAI21_X1 i_0_81 (.ZN (n_0_16), .A (n_0_90), .B1 (n_0_14), .B2 (n_0_15));
INV_X1 i_0_80 (.ZN (n_0_15), .A (n_0_94));
AOI21_X1 i_0_79 (.ZN (n_0_14), .A (n_0_13), .B1 (n_0_12), .B2 (n_0_95));
INV_X1 i_0_78 (.ZN (n_0_13), .A (n_0_98));
OAI21_X1 i_0_76 (.ZN (n_0_12), .A (n_0_11), .B1 (n_0_10), .B2 (n_0_76));
INV_X1 i_0_75 (.ZN (n_0_11), .A (n_0_97));
AOI21_X1 i_0_73 (.ZN (n_0_10), .A (n_0_227), .B1 (n_0_9), .B2 (n_0_65));
AOI21_X1 i_0_72 (.ZN (n_0_9), .A (n_0_66), .B1 (n_0_293), .B2 (n_0_8));
INV_X1 i_0_70 (.ZN (n_0_8), .A (n_0_77));
OAI21_X1 i_0_69 (.ZN (n_0_146), .A (n_0_113), .B1 (n_0_6), .B2 (n_0_7));
INV_X1 i_0_68 (.ZN (n_0_7), .A (n_0_27));
AOI21_X1 i_0_67 (.ZN (n_0_6), .A (n_0_262), .B1 (n_0_5), .B2 (n_0_263));
NAND3_X1 i_0_65 (.ZN (n_0_5), .A1 (n_0_244), .A2 (n_0_102), .A3 (n_0_110));
OAI21_X1 i_0_64 (.ZN (n_0_171), .A (n_0_4), .B1 (n_0_3), .B2 (n_0_182));
INV_X1 i_0_63 (.ZN (n_0_4), .A (n_0_139));
AOI21_X1 i_0_62 (.ZN (n_0_3), .A (n_0_2), .B1 (n_0_1), .B2 (n_0_180));
INV_X1 i_0_61 (.ZN (n_0_2), .A (n_0_138));
OAI22_X1 i_0_60 (.ZN (n_0_1), .A1 (n_0_0), .A2 (n_0_183), .B1 (i_add2[23]), .B2 (i_add1[23]));
NAND2_X1 i_0_59 (.ZN (n_0_0), .A1 (n_0_389), .A2 (n_0_189));
NAND4_X1 i_0_58 (.ZN (n_0_389), .A1 (n_0_385), .A2 (n_0_192), .A3 (n_0_144), .A4 (n_0_140));
OAI21_X1 i_0_57 (.ZN (n_0_181), .A (n_0_194), .B1 (n_0_387), .B2 (n_0_388));
INV_X1 i_0_56 (.ZN (n_0_388), .A (n_0_41));
AOI21_X1 i_0_55 (.ZN (n_0_387), .A (n_0_145), .B1 (n_0_386), .B2 (n_0_168));
NAND2_X1 i_0_54 (.ZN (n_0_386), .A1 (n_0_385), .A2 (n_0_143));
NOR2_X1 i_0_53 (.ZN (n_0_385), .A1 (n_0_384), .A2 (n_0_147));
NOR3_X1 i_0_52 (.ZN (n_0_384), .A1 (n_0_195), .A2 (n_0_184), .A3 (n_0_174));
OAI21_X1 i_0_51 (.ZN (n_0_51), .A (n_0_300), .B1 (n_0_21), .B2 (n_0_81));
AOI21_X1 i_0_50 (.ZN (n_0_301), .A (n_0_295), .B1 (n_0_299), .B2 (n_0_300));
NAND2_X1 i_0_46 (.ZN (n_0_300), .A1 (i_add1[42]), .A2 (i_add2[42]));
OAI21_X1 i_0_45 (.ZN (n_0_299), .A (n_0_80), .B1 (n_0_294), .B2 (n_0_298));
INV_X1 i_0_44 (.ZN (n_0_298), .A (n_0_21));
INV_X1 i_0_43 (.ZN (n_0_295), .A (n_0_82));
AND2_X1 i_0_42 (.ZN (n_0_294), .A1 (n_0_293), .A2 (n_0_83));
AND3_X1 i_0_41 (.ZN (n_0_293), .A1 (n_0_124), .A2 (n_0_84), .A3 (n_0_99));
AOI22_X1 i_0_40 (.ZN (n_0_50), .A1 (n_0_264), .A2 (n_0_113), .B1 (i_add1[36]), .B2 (i_add2[36]));
OAI21_X1 i_0_39 (.ZN (n_0_264), .A (n_0_27), .B1 (n_0_262), .B2 (n_0_263));
NAND2_X1 i_0_38 (.ZN (n_0_263), .A1 (i_add1[34]), .A2 (i_add2[34]));
INV_X1 i_0_37 (.ZN (n_0_262), .A (n_0_115));
AOI21_X1 i_0_35 (.ZN (n_0_261), .A (n_0_259), .B1 (n_0_326), .B2 (n_0_156));
INV_X1 i_0_34 (.ZN (n_0_259), .A (n_0_107));
NAND2_X1 i_0_33 (.ZN (n_0_49), .A1 (n_0_237), .A2 (n_0_122));
OAI21_X1 i_0_32 (.ZN (n_0_237), .A (n_0_232), .B1 (n_0_35), .B2 (n_0_120));
AOI21_X1 i_0_31 (.ZN (n_0_233), .A (n_0_202), .B1 (n_0_231), .B2 (n_0_232));
NAND2_X1 i_0_30 (.ZN (n_0_232), .A1 (i_add1[28]), .A2 (i_add2[28]));
OAI21_X1 i_0_29 (.ZN (n_0_231), .A (n_0_119), .B1 (n_0_201), .B2 (n_0_230));
INV_X1 i_0_28 (.ZN (n_0_230), .A (n_0_35));
INV_X1 i_0_27 (.ZN (n_0_202), .A (n_0_122));
AND2_X1 i_0_25 (.ZN (n_0_201), .A1 (n_0_246), .A2 (n_0_123));
OAI21_X1 i_0_188 (.ZN (n_0_48), .A (n_0_41), .B1 (n_0_145), .B2 (n_0_168));
NAND2_X1 i_0_24 (.ZN (n_0_168), .A1 (i_add1[20]), .A2 (i_add2[20]));
NAND2_X1 i_0_22 (.ZN (n_0_47), .A1 (n_0_157), .A2 (n_0_175));
OAI21_X1 i_0_21 (.ZN (n_0_157), .A (n_0_255), .B1 (n_0_256), .B2 (n_0_155));
INV_X1 i_0_20 (.ZN (n_0_155), .A (n_0_177));
INV_X1 i_0_176 (.ZN (n_0_46), .A (n_0_178));
INV_X1 i_0_166 (.ZN (n_0_45), .A (n_0_336));
INV_X1 i_0_159 (.ZN (n_0_44), .A (n_0_369));
INV_X1 i_0_97 (.ZN (w_G), .A (n_0_381));
NOR2_X1 i_0_94 (.ZN (n_23), .A1 (n_0_377), .A2 (n_0_376));
OR2_X1 i_0_91 (.ZN (n_0_42), .A1 (i_add2[4]), .A2 (i_add1[4]));
NOR2_X1 i_0_89 (.ZN (n_22), .A1 (n_0_225), .A2 (n_0_234));
NOR2_X1 i_0_19 (.ZN (n_21), .A1 (n_0_367), .A2 (n_0_372));
NOR2_X1 i_0_77 (.ZN (n_20), .A1 (n_0_363), .A2 (n_0_340));
NOR2_X1 i_0_74 (.ZN (n_19), .A1 (n_0_352), .A2 (n_0_358));
NOR2_X1 i_0_71 (.ZN (n_18), .A1 (n_0_349), .A2 (n_0_333));
INV_X1 i_0_66 (.ZN (n_17), .A (n_0_252));
INV_X1 i_0_18 (.ZN (n_16), .A (n_0_386));
NAND2_X1 i_0_17 (.ZN (n_0_41), .A1 (i_add2[21]), .A2 (i_add1[21]));
INV_X1 i_0_16 (.ZN (n_15), .A (n_0_181));
INV_X1 i_0_15 (.ZN (n_14), .A (n_0_1));
INV_X1 i_0_14 (.ZN (n_13), .A (n_0_171));
NAND2_X1 i_0_13 (.ZN (n_0_35), .A1 (i_add2[27]), .A2 (i_add1[27]));
INV_X1 i_0_12 (.ZN (n_12), .A (n_0_231));
NAND2_X1 i_0_49 (.ZN (n_0_40), .A1 (i_add2[29]), .A2 (i_add1[29]));
INV_X1 i_0_48 (.ZN (n_11), .A (n_0_245));
OR2_X1 i_0_47 (.ZN (n_0_39), .A1 (i_add2[30]), .A2 (i_add1[30]));
INV_X1 i_0_11 (.ZN (n_10), .A (n_0_5));
NAND2_X1 i_0_10 (.ZN (n_0_27), .A1 (i_add2[35]), .A2 (i_add1[35]));
INV_X1 i_0_9 (.ZN (n_9), .A (n_0_146));
INV_X1 i_0_36 (.ZN (n_8), .A (n_0_241));
NAND2_X1 i_0_8 (.ZN (n_0_21), .A1 (i_add2[41]), .A2 (i_add1[41]));
INV_X1 i_0_7 (.ZN (n_7), .A (n_0_299));
INV_X1 i_0_6 (.ZN (n_6), .A (n_0_9));
OR2_X1 i_0_26 (.ZN (n_0_38), .A1 (i_add2[44]), .A2 (i_add1[44]));
INV_X1 i_0_5 (.ZN (n_5), .A (n_0_12));
INV_X1 i_0_4 (.ZN (n_4), .A (n_0_16));
INV_X1 i_0_3 (.ZN (n_3), .A (n_0_111));
INV_X1 i_0_2 (.ZN (n_2), .A (n_0_54));
INV_X1 i_0_1 (.ZN (n_1), .A (n_0_101));
INV_X1 i_0_0 (.ZN (n_0), .A (n_0_96));
full_adder genblk1_63_full_adder_inst (.o_sum (o_result[63]), .i_bit1 (i_add1[63])
    , .i_bit2 (i_add2[63]), .i_carry (n_46));
full_adder__0_465 genblk1_62_full_adder_inst (.o_sum (o_result[62]), .i_bit1 (i_add1[62])
    , .i_bit2 (i_add2[62]), .i_carry (n_47));
full_adder__0_461 genblk1_61_full_adder_inst (.o_sum (o_result[61]), .i_bit1 (i_add1[61])
    , .i_bit2 (i_add2[61]), .i_carry (n_0_319));
full_adder__0_457 genblk1_60_full_adder_inst (.o_sum (o_result[60]), .i_bit1 (i_add1[60])
    , .i_bit2 (i_add2[60]), .i_carry (n_48));
full_adder__0_453 genblk1_59_full_adder_inst (.o_sum (o_result[59]), .i_bit1 (i_add1[59])
    , .i_bit2 (i_add2[59]), .i_carry (n_0_323));
full_adder__0_449 genblk1_58_full_adder_inst (.o_sum (o_result[58]), .i_bit1 (i_add1[58])
    , .i_bit2 (i_add2[58]), .i_carry (n_49));
full_adder__0_445 genblk1_57_full_adder_inst (.o_sum (o_result[57]), .i_bit1 (i_add1[57])
    , .i_bit2 (i_add2[57]), .i_carry (n_42));
full_adder__0_441 genblk1_56_full_adder_inst (.o_sum (o_result[56]), .i_bit1 (i_add1[56])
    , .i_bit2 (i_add2[56]), .i_carry (n_0));
full_adder__0_437 genblk1_55_full_adder_inst (.o_sum (o_result[55]), .i_bit1 (i_add1[55])
    , .i_bit2 (i_add2[55]), .i_carry (n_0_22));
full_adder__0_433 genblk1_54_full_adder_inst (.o_sum (o_result[54]), .i_bit1 (i_add1[54])
    , .i_bit2 (i_add2[54]), .i_carry (n_1));
full_adder__0_429 genblk1_53_full_adder_inst (.o_sum (o_result[53]), .i_bit1 (i_add1[53])
    , .i_bit2 (i_add2[53]), .i_carry (n_0_52));
full_adder__0_425 genblk1_52_full_adder_inst (.o_sum (o_result[52]), .i_bit1 (i_add1[52])
    , .i_bit2 (i_add2[52]), .i_carry (n_2));
full_adder__0_421 genblk1_51_full_adder_inst (.o_sum (o_result[51]), .i_bit1 (i_add1[51])
    , .i_bit2 (i_add2[51]), .i_carry (n_0_57));
full_adder__0_417 genblk1_50_full_adder_inst (.o_sum (o_result[50]), .i_bit1 (i_add1[50])
    , .i_bit2 (i_add2[50]), .i_carry (n_3));
full_adder__0_413 genblk1_49_full_adder_inst (.o_sum (o_result[49]), .i_bit1 (i_add1[49])
    , .i_bit2 (i_add2[49]), .i_carry (n_0_17));
full_adder__0_409 genblk1_48_full_adder_inst (.o_sum (o_result[48]), .i_bit1 (i_add1[48])
    , .i_bit2 (i_add2[48]), .i_carry (n_4));
full_adder__0_405 genblk1_47_full_adder_inst (.o_sum (o_result[47]), .i_bit1 (i_add1[47])
    , .i_bit2 (i_add2[47]), .i_carry (n_0_14));
full_adder__0_401 genblk1_46_full_adder_inst (.o_sum (o_result[46]), .i_bit1 (i_add1[46])
    , .i_bit2 (i_add2[46]), .i_carry (n_5));
full_adder__0_397 genblk1_45_full_adder_inst (.o_sum (o_result[45]), .i_bit1 (i_add1[45])
    , .i_bit2 (i_add2[45]), .i_carry (n_0_10));
full_adder__0_393 genblk1_44_full_adder_inst (.o_sum (o_result[44]), .i_bit1 (i_add1[44])
    , .i_bit2 (i_add2[44]), .i_carry (n_6));
full_adder__0_389 genblk1_43_full_adder_inst (.o_sum (o_result[43]), .i_bit1 (i_add1[43])
    , .i_bit2 (i_add2[43]), .i_carry (n_0_301));
full_adder__0_385 genblk1_42_full_adder_inst (.o_sum (o_result[42]), .i_bit1 (i_add1[42])
    , .i_bit2 (i_add2[42]), .i_carry (n_7));
full_adder__0_381 genblk1_41_full_adder_inst (.o_sum (o_result[41]), .i_bit1 (i_add1[41])
    , .i_bit2 (i_add2[41]), .i_carry (n_0_294));
full_adder__0_377 genblk1_40_full_adder_inst (.o_sum (o_result[40]), .i_bit1 (i_add1[40])
    , .i_bit2 (i_add2[40]), .i_carry (n_50));
full_adder__0_373 genblk1_39_full_adder_inst (.o_sum (o_result[39]), .i_bit1 (i_add1[39])
    , .i_bit2 (i_add2[39]), .i_carry (n_0_240));
full_adder__0_369 genblk1_38_full_adder_inst (.o_sum (o_result[38]), .i_bit1 (i_add1[38])
    , .i_bit2 (i_add2[38]), .i_carry (n_8));
full_adder__0_365 genblk1_37_full_adder_inst (.o_sum (o_result[37]), .i_bit1 (i_add1[37])
    , .i_bit2 (i_add2[37]), .i_carry (n_0_242));
full_adder__0_361 genblk1_36_full_adder_inst (.o_sum (o_result[36]), .i_bit1 (i_add1[36])
    , .i_bit2 (i_add2[36]), .i_carry (n_9));
full_adder__0_357 genblk1_35_full_adder_inst (.o_sum (o_result[35]), .i_bit1 (i_add1[35])
    , .i_bit2 (i_add2[35]), .i_carry (n_0_6));
full_adder__0_353 genblk1_34_full_adder_inst (.o_sum (o_result[34]), .i_bit1 (i_add1[34])
    , .i_bit2 (i_add2[34]), .i_carry (n_10));
full_adder__0_349 genblk1_33_full_adder_inst (.o_sum (o_result[33]), .i_bit1 (i_add1[33])
    , .i_bit2 (i_add2[33]), .i_carry (n_0_261));
full_adder__0_345 genblk1_32_full_adder_inst (.o_sum (o_result[32]), .i_bit1 (i_add1[32])
    , .i_bit2 (i_add2[32]), .i_carry (n_51));
full_adder__0_341 genblk1_31_full_adder_inst (.o_sum (o_result[31]), .i_bit1 (i_add1[31])
    , .i_bit2 (i_add2[31]), .i_carry (n_0_328));
full_adder__0_337 genblk1_30_full_adder_inst (.o_sum (o_result[30]), .i_bit1 (i_add1[30])
    , .i_bit2 (i_add2[30]), .i_carry (n_11));
full_adder__0_333 genblk1_29_full_adder_inst (.o_sum (o_result[29]), .i_bit1 (i_add1[29])
    , .i_bit2 (i_add2[29]), .i_carry (n_0_233));
full_adder__0_329 genblk1_28_full_adder_inst (.o_sum (o_result[28]), .i_bit1 (i_add1[28])
    , .i_bit2 (i_add2[28]), .i_carry (n_12));
full_adder__0_325 genblk1_27_full_adder_inst (.o_sum (o_result[27]), .i_bit1 (i_add1[27])
    , .i_bit2 (i_add2[27]), .i_carry (n_0_201));
full_adder__0_321 genblk1_26_full_adder_inst (.o_sum (o_result[26]), .i_bit1 (i_add1[26])
    , .i_bit2 (i_add2[26]), .i_carry (n_13));
full_adder__0_317 genblk1_25_full_adder_inst (.o_sum (o_result[25]), .i_bit1 (i_add1[25])
    , .i_bit2 (i_add2[25]), .i_carry (n_0_3));
full_adder__0_313 genblk1_24_full_adder_inst (.o_sum (o_result[24]), .i_bit1 (i_add1[24])
    , .i_bit2 (i_add2[24]), .i_carry (n_14));
full_adder__0_309 genblk1_23_full_adder_inst (.o_sum (o_result[23]), .i_bit1 (i_add1[23])
    , .i_bit2 (i_add2[23]), .i_carry (n_0_0));
full_adder__0_305 genblk1_22_full_adder_inst (.o_sum (o_result[22]), .i_bit1 (i_add1[22])
    , .i_bit2 (i_add2[22]), .i_carry (n_15));
full_adder__0_301 genblk1_21_full_adder_inst (.o_sum (o_result[21]), .i_bit1 (i_add1[21])
    , .i_bit2 (i_add2[21]), .i_carry (n_0_387));
full_adder__0_297 genblk1_20_full_adder_inst (.o_sum (o_result[20]), .i_bit1 (i_add1[20])
    , .i_bit2 (i_add2[20]), .i_carry (n_16));
full_adder__0_293 genblk1_19_full_adder_inst (.o_sum (o_result[19]), .i_bit1 (i_add1[19])
    , .i_bit2 (i_add2[19]), .i_carry (n_0_251));
full_adder__0_289 genblk1_18_full_adder_inst (.o_sum (o_result[18]), .i_bit1 (i_add1[18])
    , .i_bit2 (i_add2[18]), .i_carry (n_17));
full_adder__0_285 genblk1_17_full_adder_inst (.o_sum (o_result[17]), .i_bit1 (i_add1[17])
    , .i_bit2 (i_add2[17]), .i_carry (n_52));
full_adder__0_281 genblk1_16_full_adder_inst (.o_sum (o_result[16]), .i_bit1 (i_add1[16])
    , .i_bit2 (i_add2[16]), .i_carry (n_53));
full_adder__0_277 genblk1_15_full_adder_inst (.o_sum (o_result[15]), .i_bit1 (i_add1[15])
    , .i_bit2 (i_add2[15]), .i_carry (n_18));
full_adder__0_273 genblk1_14_full_adder_inst (.o_sum (o_result[14]), .i_bit1 (i_add1[14])
    , .i_bit2 (i_add2[14]), .i_carry (n_54));
full_adder__0_269 genblk1_13_full_adder_inst (.o_sum (o_result[13]), .i_bit1 (i_add1[13])
    , .i_bit2 (i_add2[13]), .i_carry (n_19));
full_adder__0_265 genblk1_12_full_adder_inst (.o_sum (o_result[12]), .i_bit1 (i_add1[12])
    , .i_bit2 (i_add2[12]), .i_carry (n_55));
full_adder__0_261 genblk1_11_full_adder_inst (.o_sum (o_result[11]), .i_bit1 (i_add1[11])
    , .i_bit2 (i_add2[11]), .i_carry (n_20));
full_adder__0_257 genblk1_10_full_adder_inst (.o_sum (o_result[10]), .i_bit1 (i_add1[10])
    , .i_bit2 (i_add2[10]), .i_carry (n_56));
full_adder__0_253 genblk1_9_full_adder_inst (.o_sum (o_result[9]), .i_bit1 (i_add1[9])
    , .i_bit2 (i_add2[9]), .i_carry (n_57));
full_adder__0_249 genblk1_8_full_adder_inst (.o_sum (o_result[8]), .i_bit1 (i_add1[8])
    , .i_bit2 (i_add2[8]), .i_carry (n_58));
full_adder__0_245 genblk1_7_full_adder_inst (.o_sum (o_result[7]), .i_bit1 (i_add1[7])
    , .i_bit2 (i_add2[7]), .i_carry (n_21));
full_adder__0_241 genblk1_6_full_adder_inst (.o_sum (o_result[6]), .i_bit1 (i_add1[6])
    , .i_bit2 (i_add2[6]), .i_carry (n_59));
full_adder__0_237 genblk1_5_full_adder_inst (.o_sum (o_result[5]), .i_bit1 (i_add1[5])
    , .i_bit2 (i_add2[5]), .i_carry (n_22));
full_adder__0_233 genblk1_4_full_adder_inst (.o_sum (o_result[4]), .i_bit1 (i_add1[4])
    , .i_bit2 (i_add2[4]), .i_carry (n_60));
full_adder__0_229 genblk1_3_full_adder_inst (.o_sum (o_result[3]), .i_bit1 (i_add1[3])
    , .i_bit2 (i_add2[3]), .i_carry (n_23));
full_adder__0_225 genblk1_2_full_adder_inst (.o_sum (o_result[2]), .i_bit1 (i_add1[2])
    , .i_bit2 (i_add2[2]), .i_carry (n_61));
full_adder__0_221 genblk1_1_full_adder_inst (.o_sum (o_result[1]), .i_bit1 (i_add1[1])
    , .i_bit2 (i_add2[1]), .i_carry (w_G));
full_adder__0_217 genblk1_0_full_adder_inst (.o_sum (o_result[0]), .i_bit1 (i_add1[0])
    , .i_bit2 (i_add2[0]));

endmodule //carry_lookahead_adder

module regFile (clk__CTS_1_PP_1, read_data, read_data2, write_en, write_data, write_data2, 
    clk);

output [31:0] read_data2;
output [31:0] read_data;
input clk;
input [31:0] write_data2;
input [31:0] write_data;
input write_en;
input clk__CTS_1_PP_1;
wire CTS_n_tid0_5;
wire CTS_n_tid0_6;


CLKGATETST_X8 clk_gate_my_reg2_reg (.GCK (CTS_n_tid0_6), .CK (clk__CTS_1_PP_1), .E (write_en), .SE (1'b0 ));
DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid0_5), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid0_5), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid0_5), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid0_5), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid0_5), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid0_5), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid0_5), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid0_5), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid0_5), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid0_5), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid0_5), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid0_5), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid0_5), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid0_5), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid0_5), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid0_5), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid0_5), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid0_5), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid0_5), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid0_5), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid0_5), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid0_5), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid0_5), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid0_5), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid0_5), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid0_5), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid0_5), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid0_5), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid0_5), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid0_5), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid0_5), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid0_5), .D (write_data[31]));
DFF_X1 \my_reg2_reg[0]  (.Q (read_data2[0]), .CK (CTS_n_tid0_5), .D (write_data2[0]));
DFF_X1 \my_reg2_reg[1]  (.Q (read_data2[1]), .CK (CTS_n_tid0_5), .D (write_data2[1]));
DFF_X1 \my_reg2_reg[2]  (.Q (read_data2[2]), .CK (CTS_n_tid0_5), .D (write_data2[2]));
DFF_X1 \my_reg2_reg[3]  (.Q (read_data2[3]), .CK (CTS_n_tid0_5), .D (write_data2[3]));
DFF_X1 \my_reg2_reg[4]  (.Q (read_data2[4]), .CK (CTS_n_tid0_5), .D (write_data2[4]));
DFF_X1 \my_reg2_reg[5]  (.Q (read_data2[5]), .CK (CTS_n_tid0_5), .D (write_data2[5]));
DFF_X1 \my_reg2_reg[6]  (.Q (read_data2[6]), .CK (CTS_n_tid0_5), .D (write_data2[6]));
DFF_X1 \my_reg2_reg[7]  (.Q (read_data2[7]), .CK (CTS_n_tid0_5), .D (write_data2[7]));
DFF_X1 \my_reg2_reg[8]  (.Q (read_data2[8]), .CK (CTS_n_tid0_5), .D (write_data2[8]));
DFF_X1 \my_reg2_reg[9]  (.Q (read_data2[9]), .CK (CTS_n_tid0_5), .D (write_data2[9]));
DFF_X1 \my_reg2_reg[10]  (.Q (read_data2[10]), .CK (CTS_n_tid0_5), .D (write_data2[10]));
DFF_X1 \my_reg2_reg[11]  (.Q (read_data2[11]), .CK (CTS_n_tid0_5), .D (write_data2[11]));
DFF_X1 \my_reg2_reg[12]  (.Q (read_data2[12]), .CK (CTS_n_tid0_5), .D (write_data2[12]));
DFF_X1 \my_reg2_reg[13]  (.Q (read_data2[13]), .CK (CTS_n_tid0_5), .D (write_data2[13]));
DFF_X1 \my_reg2_reg[14]  (.Q (read_data2[14]), .CK (CTS_n_tid0_5), .D (write_data2[14]));
DFF_X1 \my_reg2_reg[15]  (.Q (read_data2[15]), .CK (CTS_n_tid0_5), .D (write_data2[15]));
DFF_X1 \my_reg2_reg[16]  (.Q (read_data2[16]), .CK (CTS_n_tid0_5), .D (write_data2[16]));
DFF_X1 \my_reg2_reg[17]  (.Q (read_data2[17]), .CK (CTS_n_tid0_5), .D (write_data2[17]));
DFF_X1 \my_reg2_reg[18]  (.Q (read_data2[18]), .CK (CTS_n_tid0_5), .D (write_data2[18]));
DFF_X1 \my_reg2_reg[19]  (.Q (read_data2[19]), .CK (CTS_n_tid0_5), .D (write_data2[19]));
DFF_X1 \my_reg2_reg[20]  (.Q (read_data2[20]), .CK (CTS_n_tid0_5), .D (write_data2[20]));
DFF_X1 \my_reg2_reg[21]  (.Q (read_data2[21]), .CK (CTS_n_tid0_5), .D (write_data2[21]));
DFF_X1 \my_reg2_reg[22]  (.Q (read_data2[22]), .CK (CTS_n_tid0_5), .D (write_data2[22]));
DFF_X1 \my_reg2_reg[23]  (.Q (read_data2[23]), .CK (CTS_n_tid0_5), .D (write_data2[23]));
DFF_X1 \my_reg2_reg[24]  (.Q (read_data2[24]), .CK (CTS_n_tid0_5), .D (write_data2[24]));
DFF_X1 \my_reg2_reg[25]  (.Q (read_data2[25]), .CK (CTS_n_tid0_5), .D (write_data2[25]));
DFF_X1 \my_reg2_reg[26]  (.Q (read_data2[26]), .CK (CTS_n_tid0_5), .D (write_data2[26]));
DFF_X1 \my_reg2_reg[27]  (.Q (read_data2[27]), .CK (CTS_n_tid0_5), .D (write_data2[27]));
DFF_X1 \my_reg2_reg[28]  (.Q (read_data2[28]), .CK (CTS_n_tid0_5), .D (write_data2[28]));
DFF_X1 \my_reg2_reg[29]  (.Q (read_data2[29]), .CK (CTS_n_tid0_5), .D (write_data2[29]));
DFF_X1 \my_reg2_reg[30]  (.Q (read_data2[30]), .CK (CTS_n_tid0_5), .D (write_data2[30]));
DFF_X1 \my_reg2_reg[31]  (.Q (read_data2[31]), .CK (CTS_n_tid0_5), .D (write_data2[31]));
CLKBUF_X3 CTS_L3_c_tid0_3 (.Z (CTS_n_tid0_5), .A (CTS_n_tid0_6));

endmodule //regFile

module Radix4 (a, b, read_data3, clk, start, start_shift, start_i);

output [63:0] read_data3;
input [31:0] a;
input [31:0] b;
input clk;
input start;
input [4:0] start_i;
input [4:0] start_shift;
wire \read_data2[31] ;
wire \read_data2[30] ;
wire \read_data2[29] ;
wire \read_data2[28] ;
wire \read_data2[27] ;
wire \read_data2[26] ;
wire \read_data2[25] ;
wire \read_data2[24] ;
wire \read_data2[23] ;
wire \read_data2[22] ;
wire \read_data2[21] ;
wire \read_data2[20] ;
wire \read_data2[19] ;
wire \read_data2[18] ;
wire \read_data2[17] ;
wire \read_data2[16] ;
wire \read_data2[15] ;
wire \read_data2[14] ;
wire \read_data2[13] ;
wire \read_data2[12] ;
wire \read_data2[11] ;
wire \read_data2[10] ;
wire \read_data2[9] ;
wire \read_data2[8] ;
wire \read_data2[7] ;
wire \read_data2[6] ;
wire \read_data2[5] ;
wire \read_data2[4] ;
wire \read_data2[3] ;
wire \read_data2[2] ;
wire \read_data2[1] ;
wire \read_data2[0] ;
wire \read_data[31] ;
wire \read_data[30] ;
wire \read_data[29] ;
wire \read_data[28] ;
wire \read_data[27] ;
wire \read_data[26] ;
wire \read_data[25] ;
wire \read_data[24] ;
wire \read_data[23] ;
wire \read_data[22] ;
wire \read_data[21] ;
wire \read_data[20] ;
wire \read_data[19] ;
wire \read_data[18] ;
wire \read_data[17] ;
wire \read_data[16] ;
wire \read_data[15] ;
wire \read_data[14] ;
wire \read_data[13] ;
wire \read_data[12] ;
wire \read_data[11] ;
wire \read_data[10] ;
wire \read_data[9] ;
wire \read_data[8] ;
wire \read_data[7] ;
wire \read_data[6] ;
wire \read_data[5] ;
wire \read_data[4] ;
wire \read_data[3] ;
wire \read_data[2] ;
wire \read_data[1] ;
wire \read_data[0] ;
wire \res[63] ;
wire \res[62] ;
wire \res[61] ;
wire \res[60] ;
wire \res[59] ;
wire \res[58] ;
wire \res[57] ;
wire \res[56] ;
wire \res[55] ;
wire \res[54] ;
wire \res[53] ;
wire \res[52] ;
wire \res[51] ;
wire \res[50] ;
wire \res[49] ;
wire \res[48] ;
wire \res[47] ;
wire \res[46] ;
wire \res[45] ;
wire \res[44] ;
wire \res[43] ;
wire \res[42] ;
wire \res[41] ;
wire \res[40] ;
wire \res[39] ;
wire \res[38] ;
wire \res[37] ;
wire \res[36] ;
wire \res[35] ;
wire \res[34] ;
wire \res[33] ;
wire \res[32] ;
wire \res[31] ;
wire \res[30] ;
wire \res[29] ;
wire \res[28] ;
wire \res[27] ;
wire \res[26] ;
wire \res[25] ;
wire \res[24] ;
wire \res[23] ;
wire \res[22] ;
wire \res[21] ;
wire \res[20] ;
wire \res[19] ;
wire \res[18] ;
wire \res[17] ;
wire \res[16] ;
wire \res[15] ;
wire \res[14] ;
wire \res[13] ;
wire \res[12] ;
wire \res[11] ;
wire \res[10] ;
wire \res[9] ;
wire \res[8] ;
wire \res[7] ;
wire \res[6] ;
wire \res[5] ;
wire \res[4] ;
wire \res[3] ;
wire \res[2] ;
wire \res[1] ;
wire \res[0] ;
wire \sum[63] ;
wire \sum[62] ;
wire \sum[61] ;
wire \sum[60] ;
wire \sum[59] ;
wire \sum[58] ;
wire \sum[57] ;
wire \sum[56] ;
wire \sum[55] ;
wire \sum[54] ;
wire \sum[53] ;
wire \sum[52] ;
wire \sum[51] ;
wire \sum[50] ;
wire \sum[49] ;
wire \sum[48] ;
wire \sum[47] ;
wire \sum[46] ;
wire \sum[45] ;
wire \sum[44] ;
wire \sum[43] ;
wire \sum[42] ;
wire \sum[41] ;
wire \sum[40] ;
wire \sum[39] ;
wire \sum[38] ;
wire \sum[37] ;
wire \sum[36] ;
wire \sum[35] ;
wire \sum[34] ;
wire \sum[33] ;
wire \sum[32] ;
wire \sum[31] ;
wire \sum[30] ;
wire \sum[29] ;
wire \sum[28] ;
wire \sum[27] ;
wire \sum[26] ;
wire \sum[25] ;
wire \sum[24] ;
wire \sum[23] ;
wire \sum[22] ;
wire \sum[21] ;
wire \sum[20] ;
wire \sum[19] ;
wire \sum[18] ;
wire \sum[17] ;
wire \sum[16] ;
wire \sum[15] ;
wire \sum[14] ;
wire \sum[13] ;
wire \sum[12] ;
wire \sum[11] ;
wire \sum[10] ;
wire \sum[9] ;
wire \sum[8] ;
wire \sum[7] ;
wire \sum[6] ;
wire \sum[5] ;
wire \sum[4] ;
wire \sum[3] ;
wire \sum[2] ;
wire \sum[1] ;
wire \sum[0] ;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_0_0;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_0_1;
wire n_0_126;
wire n_0_0_2;
wire n_0_127;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_128;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_129;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_130;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_131;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire n_0_0_60;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_0_65;
wire n_0_0_66;
wire n_0_0_67;
wire n_0_0_68;
wire n_0_0_69;
wire n_0_0_70;
wire n_0_0_71;
wire n_0_0_72;
wire n_0_0_73;
wire n_0_0_74;
wire n_0_0_75;
wire n_0_176;
wire n_0_0_76;
wire n_0_0_77;
wire n_0_0_78;
wire n_0_0_79;
wire n_0_0_80;
wire n_0_0_81;
wire n_0_0_82;
wire n_0_0_83;
wire n_0_0_84;
wire n_0_0_85;
wire n_0_0_86;
wire n_0_0_87;
wire n_0_0_88;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_93;
wire n_0_177;
wire n_0_0_94;
wire n_0_0_95;
wire n_0_0_96;
wire n_0_0_97;
wire n_0_0_98;
wire n_0_0_99;
wire n_0_0_100;
wire n_0_0_101;
wire n_0_0_102;
wire n_0_0_103;
wire n_0_178;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_179;
wire n_0_0_110;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_0_113;
wire n_0_0_114;
wire n_0_0_115;
wire n_0_0_116;
wire n_0_0_117;
wire n_0_180;
wire n_0_0_118;
wire n_0_0_119;
wire n_0_0_120;
wire n_0_0_121;
wire n_0_0_122;
wire n_0_0_123;
wire n_0_181;
wire n_0_0_124;
wire n_0_0_125;
wire n_0_0_126;
wire n_0_0_127;
wire n_0_0_128;
wire n_0_0_129;
wire n_0_0_130;
wire n_0_182;
wire n_0_0_131;
wire n_0_0_132;
wire n_0_0_133;
wire n_0_0_134;
wire n_0_0_135;
wire n_0_0_136;
wire n_0_0_137;
wire n_0_183;
wire n_0_0_138;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_144;
wire n_0_0_145;
wire n_0_0_146;
wire n_0_184;
wire n_0_0_147;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_185;
wire n_0_0_153;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_186;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_187;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_188;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_189;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_190;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_0_188;
wire n_0_191;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_192;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_0_207;
wire n_0_193;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_194;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_195;
wire n_0_0_224;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_196;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_197;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_198;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_0_248;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_199;
wire n_0_0_253;
wire n_0_0_254;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_200;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_201;
wire n_0_0_271;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_132;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_133;
wire n_0_0_289;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_134;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_0_299;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_135;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_136;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_137;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_138;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_139;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_0_339;
wire n_0_140;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_141;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_0_347;
wire n_0_142;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_143;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_0_355;
wire n_0_144;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire n_0_145;
wire n_0_0_360;
wire n_0_0_361;
wire n_0_0_362;
wire n_0_0_363;
wire n_0_0_364;
wire n_0_0_365;
wire n_0_146;
wire n_0_0_366;
wire n_0_0_367;
wire n_0_0_368;
wire n_0_147;
wire n_0_0_369;
wire n_0_0_370;
wire n_0_0_371;
wire n_0_148;
wire n_0_0_372;
wire n_0_0_373;
wire n_0_0_374;
wire n_0_149;
wire n_0_0_375;
wire n_0_0_376;
wire n_0_0_377;
wire n_0_0_378;
wire n_0_150;
wire n_0_0_379;
wire n_0_0_380;
wire n_0_0_381;
wire n_0_0_382;
wire n_0_151;
wire n_0_0_383;
wire n_0_0_384;
wire n_0_0_385;
wire n_0_0_386;
wire n_0_152;
wire n_0_0_387;
wire n_0_0_388;
wire n_0_0_389;
wire n_0_0_390;
wire n_0_153;
wire n_0_0_391;
wire n_0_0_392;
wire n_0_0_393;
wire n_0_0_394;
wire n_0_154;
wire n_0_0_395;
wire n_0_0_396;
wire n_0_0_397;
wire n_0_155;
wire n_0_0_398;
wire n_0_0_399;
wire n_0_0_400;
wire n_0_156;
wire n_0_0_401;
wire n_0_0_402;
wire n_0_0_403;
wire n_0_157;
wire n_0_0_404;
wire n_0_0_405;
wire n_0_0_406;
wire n_0_0_407;
wire n_0_158;
wire n_0_0_408;
wire n_0_0_409;
wire n_0_0_410;
wire n_0_0_411;
wire n_0_0_412;
wire n_0_159;
wire n_0_0_413;
wire n_0_0_414;
wire n_0_0_415;
wire n_0_160;
wire n_0_0_416;
wire n_0_0_417;
wire n_0_0_418;
wire n_0_0_419;
wire n_0_0_420;
wire n_0_161;
wire n_0_0_421;
wire n_0_0_422;
wire n_0_0_423;
wire n_0_0_424;
wire n_0_162;
wire n_0_0_425;
wire n_0_0_426;
wire n_0_0_427;
wire n_0_0_428;
wire n_0_163;
wire n_0_0_429;
wire n_0_0_430;
wire n_0_164;
wire n_0_0_431;
wire n_0_0_432;
wire n_0_165;
wire n_0_0_433;
wire n_0_0_434;
wire n_0_0_435;
wire n_0_0_436;
wire n_0_0_437;
wire n_0_0_438;
wire n_0_0_439;
wire n_0_166;
wire n_0_0_440;
wire n_0_0_441;
wire n_0_167;
wire n_0_169;
wire n_0_0_442;
wire n_0_168;
wire n_0_0_443;
wire n_0_170;
wire n_0_0_444;
wire n_0_171;
wire n_0_0_445;
wire n_0_0_446;
wire n_0_172;
wire n_0_0_447;
wire n_0_0_448;
wire n_0_173;
wire n_0_0_449;
wire n_0_0_450;
wire n_0_174;
wire write_en;
wire \c[63] ;
wire \c[62] ;
wire \c[61] ;
wire \c[60] ;
wire \c[59] ;
wire \c[58] ;
wire \c[57] ;
wire \c[56] ;
wire \c[55] ;
wire \c[54] ;
wire \c[53] ;
wire \c[52] ;
wire \c[51] ;
wire \c[50] ;
wire \c[49] ;
wire \c[48] ;
wire \c[47] ;
wire \c[46] ;
wire \c[45] ;
wire \c[44] ;
wire \c[43] ;
wire \c[42] ;
wire \c[41] ;
wire \c[40] ;
wire \c[39] ;
wire \c[38] ;
wire \c[37] ;
wire \c[36] ;
wire \c[35] ;
wire \c[34] ;
wire \c[33] ;
wire \c[32] ;
wire \c[31] ;
wire \c[30] ;
wire \c[29] ;
wire \c[28] ;
wire \c[27] ;
wire \c[26] ;
wire \c[25] ;
wire \c[24] ;
wire \c[23] ;
wire \c[22] ;
wire \c[21] ;
wire \c[20] ;
wire \c[19] ;
wire \c[18] ;
wire \c[17] ;
wire \c[16] ;
wire \c[15] ;
wire \c[14] ;
wire \c[13] ;
wire \c[12] ;
wire \c[11] ;
wire \c[10] ;
wire \c[9] ;
wire \c[8] ;
wire \c[7] ;
wire \c[6] ;
wire \c[5] ;
wire \c[4] ;
wire \c[3] ;
wire \c[2] ;
wire \c[1] ;
wire \c[0] ;
wire \shift[4] ;
wire \shift[3] ;
wire \shift[2] ;
wire \shift[1] ;
wire \shift[0] ;
wire \i[4] ;
wire \i[3] ;
wire \i[2] ;
wire \i[1] ;
wire \i[0] ;
wire n_0_175;
wire uc_0;
wire uc_1;
wire uc_2;
wire CTS_n_tid1_74;
wire hfn_ipo_n24;
wire hfn_ipo_n32;
wire drc_ipo_n33;
wire hfn_ipo_n25;
wire n_tid1_110;
wire hfn_ipo_n27;
wire CTS_n_tid1_55;
wire hfn_ipo_n31;
wire hfn_ipo_n29;
wire drc_ipo_n34;
wire CTS_n_tid1_75;


CLKGATETST_X1 clk_gate_i_reg (.GCK (n_0_175), .CK (n_tid1_110), .E (n_0_131), .SE (1'b0 ));
DFF_X1 \i_reg[0]  (.Q (\i[0] ), .CK (n_0_175), .D (n_0_126));
DFF_X1 \i_reg[1]  (.Q (\i[1] ), .CK (n_0_175), .D (n_0_127));
DFF_X1 \i_reg[2]  (.Q (\i[2] ), .CK (n_0_175), .D (n_0_128));
DFF_X1 \i_reg[3]  (.Q (\i[3] ), .CK (n_0_175), .D (n_0_129));
DFF_X1 \i_reg[4]  (.Q (\i[4] ), .CK (n_0_175), .D (n_0_130));
DFF_X1 \shift_reg[0]  (.Q (\shift[0] ), .CK (n_0_175), .D (n_0_170));
DFF_X1 \shift_reg[1]  (.Q (\shift[1] ), .CK (n_0_175), .D (n_0_171));
DFF_X1 \shift_reg[2]  (.Q (\shift[2] ), .CK (n_0_175), .D (n_0_172));
DFF_X1 \shift_reg[3]  (.Q (\shift[3] ), .CK (n_0_175), .D (n_0_173));
DFF_X1 \shift_reg[4]  (.Q (\shift[4] ), .CK (n_0_175), .D (n_0_174));
DFF_X1 \c_reg[0]  (.Q (\c[0] ), .CK (CTS_n_tid1_74), .D (n_0_0));
DFF_X1 \c_reg[1]  (.Q (\c[1] ), .CK (CTS_n_tid1_74), .D (n_0_1));
DFF_X1 \c_reg[2]  (.Q (\c[2] ), .CK (CTS_n_tid1_74), .D (n_0_2));
DFF_X1 \c_reg[3]  (.Q (\c[3] ), .CK (CTS_n_tid1_74), .D (n_0_3));
DFF_X1 \c_reg[4]  (.Q (\c[4] ), .CK (CTS_n_tid1_74), .D (n_0_4));
DFF_X1 \c_reg[5]  (.Q (\c[5] ), .CK (CTS_n_tid1_74), .D (n_0_5));
DFF_X1 \c_reg[6]  (.Q (\c[6] ), .CK (CTS_n_tid1_74), .D (n_0_6));
DFF_X1 \c_reg[7]  (.Q (\c[7] ), .CK (CTS_n_tid1_74), .D (n_0_7));
DFF_X1 \c_reg[8]  (.Q (\c[8] ), .CK (CTS_n_tid1_74), .D (n_0_8));
DFF_X1 \c_reg[9]  (.Q (\c[9] ), .CK (CTS_n_tid1_74), .D (n_0_71));
DFF_X1 \c_reg[10]  (.Q (\c[10] ), .CK (CTS_n_tid1_74), .D (n_0_72));
DFF_X1 \c_reg[11]  (.Q (\c[11] ), .CK (CTS_n_tid1_74), .D (n_0_73));
DFF_X1 \c_reg[12]  (.Q (\c[12] ), .CK (CTS_n_tid1_74), .D (n_0_74));
DFF_X1 \c_reg[13]  (.Q (\c[13] ), .CK (CTS_n_tid1_74), .D (n_0_75));
DFF_X1 \c_reg[14]  (.Q (\c[14] ), .CK (CTS_n_tid1_74), .D (n_0_76));
DFF_X1 \c_reg[15]  (.Q (\c[15] ), .CK (CTS_n_tid1_74), .D (n_0_77));
DFF_X1 \c_reg[16]  (.Q (\c[16] ), .CK (CTS_n_tid1_74), .D (n_0_78));
DFF_X1 \c_reg[17]  (.Q (\c[17] ), .CK (CTS_n_tid1_74), .D (n_0_79));
DFF_X1 \c_reg[18]  (.Q (\c[18] ), .CK (CTS_n_tid1_75), .D (n_0_80));
DFF_X1 \c_reg[19]  (.Q (\c[19] ), .CK (CTS_n_tid1_75), .D (n_0_81));
DFF_X1 \c_reg[20]  (.Q (\c[20] ), .CK (CTS_n_tid1_75), .D (n_0_82));
DFF_X1 \c_reg[21]  (.Q (\c[21] ), .CK (CTS_n_tid1_75), .D (n_0_83));
DFF_X1 \c_reg[22]  (.Q (\c[22] ), .CK (CTS_n_tid1_75), .D (n_0_84));
DFF_X1 \c_reg[23]  (.Q (\c[23] ), .CK (CTS_n_tid1_75), .D (n_0_85));
DFF_X1 \c_reg[24]  (.Q (\c[24] ), .CK (CTS_n_tid1_75), .D (n_0_86));
DFF_X1 \c_reg[25]  (.Q (\c[25] ), .CK (CTS_n_tid1_75), .D (n_0_87));
DFF_X1 \c_reg[26]  (.Q (\c[26] ), .CK (CTS_n_tid1_75), .D (n_0_88));
DFF_X1 \c_reg[27]  (.Q (\c[27] ), .CK (CTS_n_tid1_75), .D (n_0_89));
DFF_X1 \c_reg[28]  (.Q (\c[28] ), .CK (CTS_n_tid1_75), .D (n_0_90));
DFF_X1 \c_reg[29]  (.Q (\c[29] ), .CK (CTS_n_tid1_75), .D (n_0_91));
DFF_X1 \c_reg[30]  (.Q (\c[30] ), .CK (CTS_n_tid1_75), .D (n_0_92));
DFF_X1 \c_reg[31]  (.Q (\c[31] ), .CK (CTS_n_tid1_75), .D (n_0_93));
DFF_X1 \c_reg[32]  (.Q (\c[32] ), .CK (CTS_n_tid1_75), .D (n_0_94));
DFF_X1 \c_reg[33]  (.Q (\c[33] ), .CK (CTS_n_tid1_75), .D (n_0_95));
DFF_X1 \c_reg[34]  (.Q (\c[34] ), .CK (CTS_n_tid1_75), .D (n_0_96));
DFF_X1 \c_reg[35]  (.Q (\c[35] ), .CK (CTS_n_tid1_75), .D (n_0_97));
DFF_X1 \c_reg[36]  (.Q (\c[36] ), .CK (CTS_n_tid1_75), .D (n_0_98));
DFF_X1 \c_reg[37]  (.Q (\c[37] ), .CK (CTS_n_tid1_75), .D (n_0_99));
DFF_X1 \c_reg[38]  (.Q (\c[38] ), .CK (CTS_n_tid1_75), .D (n_0_100));
DFF_X1 \c_reg[39]  (.Q (\c[39] ), .CK (CTS_n_tid1_75), .D (n_0_101));
DFF_X1 \c_reg[40]  (.Q (\c[40] ), .CK (CTS_n_tid1_55), .D (n_0_102));
DFF_X1 \c_reg[41]  (.Q (\c[41] ), .CK (CTS_n_tid1_55), .D (n_0_103));
DFF_X1 \c_reg[42]  (.Q (\c[42] ), .CK (CTS_n_tid1_55), .D (n_0_104));
DFF_X1 \c_reg[43]  (.Q (\c[43] ), .CK (CTS_n_tid1_55), .D (n_0_105));
DFF_X1 \c_reg[44]  (.Q (\c[44] ), .CK (CTS_n_tid1_55), .D (n_0_106));
DFF_X1 \c_reg[45]  (.Q (\c[45] ), .CK (CTS_n_tid1_55), .D (n_0_107));
DFF_X1 \c_reg[46]  (.Q (\c[46] ), .CK (CTS_n_tid1_55), .D (n_0_108));
DFF_X1 \c_reg[47]  (.Q (\c[47] ), .CK (CTS_n_tid1_55), .D (n_0_109));
DFF_X1 \c_reg[48]  (.Q (\c[48] ), .CK (CTS_n_tid1_55), .D (n_0_110));
DFF_X1 \c_reg[49]  (.Q (\c[49] ), .CK (CTS_n_tid1_55), .D (n_0_111));
DFF_X1 \c_reg[50]  (.Q (\c[50] ), .CK (CTS_n_tid1_55), .D (n_0_112));
DFF_X1 \c_reg[51]  (.Q (\c[51] ), .CK (CTS_n_tid1_55), .D (n_0_113));
DFF_X1 \c_reg[52]  (.Q (\c[52] ), .CK (CTS_n_tid1_55), .D (n_0_114));
DFF_X1 \c_reg[53]  (.Q (\c[53] ), .CK (CTS_n_tid1_55), .D (n_0_115));
DFF_X1 \c_reg[54]  (.Q (\c[54] ), .CK (CTS_n_tid1_55), .D (n_0_116));
DFF_X1 \c_reg[55]  (.Q (\c[55] ), .CK (CTS_n_tid1_55), .D (n_0_117));
DFF_X1 \c_reg[56]  (.Q (\c[56] ), .CK (CTS_n_tid1_55), .D (n_0_118));
DFF_X1 \c_reg[57]  (.Q (\c[57] ), .CK (CTS_n_tid1_55), .D (n_0_119));
DFF_X1 \c_reg[58]  (.Q (\c[58] ), .CK (CTS_n_tid1_55), .D (n_0_120));
DFF_X1 \c_reg[59]  (.Q (\c[59] ), .CK (CTS_n_tid1_55), .D (n_0_121));
DFF_X1 \c_reg[60]  (.Q (\c[60] ), .CK (CTS_n_tid1_55), .D (n_0_122));
DFF_X1 \c_reg[61]  (.Q (\c[61] ), .CK (CTS_n_tid1_55), .D (n_0_123));
DFF_X1 \c_reg[62]  (.Q (\c[62] ), .CK (CTS_n_tid1_55), .D (n_0_124));
DFF_X1 \c_reg[63]  (.Q (\c[63] ), .CK (CTS_n_tid1_55), .D (n_0_125));
DFF_X1 write_en_reg (.Q (write_en), .CK (CTS_n_tid1_55), .D (start));
NAND2_X1 i_0_0_589 (.ZN (n_0_174), .A1 (n_0_0_449), .A2 (n_0_0_450));
NAND2_X1 i_0_0_588 (.ZN (n_0_0_450), .A1 (start), .A2 (start_shift[4]));
OAI211_X1 i_0_0_587 (.ZN (n_0_0_449), .A (n_0_0_437), .B (n_0_0_0), .C1 (\shift[4] ), .C2 (n_0_0_436));
OAI21_X1 i_0_0_586 (.ZN (n_0_173), .A (n_0_0_447), .B1 (n_0_0_448), .B2 (start));
OAI21_X1 i_0_0_585 (.ZN (n_0_0_448), .A (n_0_0_435), .B1 (drc_ipo_n34), .B2 (n_0_0_434));
NAND2_X1 i_0_0_584 (.ZN (n_0_0_447), .A1 (start_shift[3]), .A2 (start));
NAND2_X1 i_0_0_583 (.ZN (n_0_172), .A1 (n_0_0_445), .A2 (n_0_0_446));
NAND2_X1 i_0_0_582 (.ZN (n_0_0_446), .A1 (start_shift[2]), .A2 (start));
OAI211_X1 i_0_0_581 (.ZN (n_0_0_445), .A (n_0_0_433), .B (n_0_0_0), .C1 (drc_ipo_n33), .C2 (hfn_ipo_n32));
AOI22_X1 i_0_0_580 (.ZN (n_0_171), .A1 (n_0_0_444), .A2 (start), .B1 (n_0_0_0), .B2 (hfn_ipo_n32));
INV_X1 i_0_0_579 (.ZN (n_0_0_444), .A (start_shift[1]));
INV_X1 i_0_0_578 (.ZN (n_0_170), .A (n_0_0_443));
OAI22_X1 i_0_0_577 (.ZN (n_0_0_443), .A1 (n_0_0_0), .A2 (start_shift[0]), .B1 (\shift[0] ), .B2 (start));
AOI22_X1 i_0_0_576 (.ZN (n_0_168), .A1 (n_0_0_441), .A2 (\shift[0] ), .B1 (n_0_0_109), .B2 (n_0_0_442));
INV_X1 i_0_0_575 (.ZN (n_0_0_442), .A (n_0_169));
NOR2_X1 i_0_0_574 (.ZN (n_0_169), .A1 (n_0_0_321), .A2 (n_0_0_94));
OAI22_X1 i_0_0_573 (.ZN (n_0_167), .A1 (n_0_0_439), .A2 (n_0_0_109), .B1 (n_0_0_441), .B2 (n_0_0_108));
OAI21_X1 i_0_0_572 (.ZN (n_0_0_441), .A (n_0_0_438), .B1 (n_0_0_440), .B2 (n_0_0_437));
INV_X1 i_0_0_571 (.ZN (n_0_0_440), .A (n_0_0_315));
OAI22_X1 i_0_0_570 (.ZN (n_0_166), .A1 (n_0_0_432), .A2 (n_0_0_109), .B1 (n_0_0_439), .B2 (n_0_0_108));
OAI21_X1 i_0_0_569 (.ZN (n_0_0_439), .A (n_0_0_438), .B1 (n_0_0_101), .B2 (n_0_0_429));
NAND2_X1 i_0_0_568 (.ZN (n_0_0_438), .A1 (n_0_0_321), .A2 (n_0_0_437));
NAND2_X1 i_0_0_567 (.ZN (n_0_0_437), .A1 (n_0_0_436), .A2 (\shift[4] ));
INV_X1 i_0_0_566 (.ZN (n_0_0_436), .A (n_0_0_435));
NAND2_X1 i_0_0_565 (.ZN (n_0_0_435), .A1 (n_0_0_434), .A2 (drc_ipo_n34));
INV_X1 i_0_0_564 (.ZN (n_0_0_434), .A (n_0_0_433));
NAND2_X1 i_0_0_563 (.ZN (n_0_0_433), .A1 (drc_ipo_n33), .A2 (hfn_ipo_n32));
OAI22_X1 i_0_0_562 (.ZN (n_0_165), .A1 (n_0_0_430), .A2 (n_0_0_109), .B1 (n_0_0_432), .B2 (n_0_0_108));
OAI21_X1 i_0_0_561 (.ZN (n_0_0_432), .A (n_0_0_421), .B1 (n_0_0_431), .B2 (n_0_0_417));
OAI22_X1 i_0_0_560 (.ZN (n_0_0_431), .A1 (n_0_0_315), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_299));
OAI22_X1 i_0_0_559 (.ZN (n_0_164), .A1 (n_0_0_428), .A2 (n_0_0_109), .B1 (n_0_0_430), .B2 (n_0_0_108));
AOI22_X1 i_0_0_558 (.ZN (n_0_0_430), .A1 (n_0_0_423), .A2 (hfn_ipo_n32), .B1 (n_0_0_425), .B2 (n_0_0_429));
NAND2_X1 i_0_0_557 (.ZN (n_0_0_429), .A1 (n_0_0_307), .A2 (n_0_0_418));
OAI22_X1 i_0_0_556 (.ZN (n_0_163), .A1 (n_0_0_428), .A2 (n_0_0_108), .B1 (n_0_0_424), .B2 (n_0_0_109));
AOI21_X1 i_0_0_555 (.ZN (n_0_0_428), .A (n_0_0_427), .B1 (n_0_0_419), .B2 (hfn_ipo_n32));
AOI21_X1 i_0_0_554 (.ZN (n_0_0_427), .A (n_0_0_426), .B1 (n_0_0_299), .B2 (n_0_0_418));
INV_X1 i_0_0_553 (.ZN (n_0_0_426), .A (n_0_0_425));
NOR2_X1 i_0_0_552 (.ZN (n_0_0_425), .A1 (n_0_0_422), .A2 (hfn_ipo_n32));
OAI22_X1 i_0_0_551 (.ZN (n_0_162), .A1 (n_0_0_420), .A2 (n_0_0_109), .B1 (n_0_0_424), .B2 (n_0_0_108));
AOI22_X1 i_0_0_550 (.ZN (n_0_0_424), .A1 (n_0_0_414), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_423));
AOI21_X1 i_0_0_549 (.ZN (n_0_0_423), .A (n_0_0_422), .B1 (n_0_0_292), .B2 (n_0_0_418));
INV_X1 i_0_0_548 (.ZN (n_0_0_422), .A (n_0_0_421));
NAND2_X1 i_0_0_547 (.ZN (n_0_0_421), .A1 (n_0_0_321), .A2 (n_0_0_417));
OAI22_X1 i_0_0_546 (.ZN (n_0_161), .A1 (n_0_0_420), .A2 (n_0_0_108), .B1 (n_0_0_415), .B2 (n_0_0_109));
OAI22_X1 i_0_0_545 (.ZN (n_0_0_420), .A1 (n_0_0_411), .A2 (n_0_0_101), .B1 (n_0_0_419), .B2 (hfn_ipo_n32));
AOI221_X1 i_0_0_544 (.ZN (n_0_0_419), .A (n_0_0_416), .B1 (n_0_0_315), .B2 (n_0_0_404)
    , .C1 (n_0_0_283), .C2 (n_0_0_418));
INV_X1 i_0_0_543 (.ZN (n_0_0_418), .A (n_0_0_417));
NAND2_X1 i_0_0_542 (.ZN (n_0_0_417), .A1 (n_0_0_362), .A2 (drc_ipo_n33));
INV_X1 i_0_0_541 (.ZN (n_0_0_416), .A (n_0_0_391));
OAI22_X1 i_0_0_540 (.ZN (n_0_160), .A1 (n_0_0_412), .A2 (n_0_0_109), .B1 (n_0_0_415), .B2 (n_0_0_108));
AOI22_X1 i_0_0_539 (.ZN (n_0_0_415), .A1 (n_0_0_414), .A2 (n_0_0_101), .B1 (hfn_ipo_n32), .B2 (n_0_0_406));
AOI22_X1 i_0_0_538 (.ZN (n_0_0_414), .A1 (n_0_0_413), .A2 (n_0_0_410), .B1 (drc_ipo_n33), .B2 (n_0_0_398));
NAND2_X1 i_0_0_537 (.ZN (n_0_0_413), .A1 (n_0_0_383), .A2 (drc_ipo_n34));
OAI22_X1 i_0_0_536 (.ZN (n_0_159), .A1 (n_0_0_407), .A2 (n_0_0_109), .B1 (n_0_0_412), .B2 (n_0_0_108));
OAI22_X1 i_0_0_535 (.ZN (n_0_0_412), .A1 (n_0_0_402), .A2 (n_0_0_101), .B1 (n_0_0_411), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_0_534 (.ZN (n_0_0_411), .A1 (n_0_0_408), .A2 (n_0_0_410), .B1 (drc_ipo_n33), .B2 (n_0_0_395));
AOI21_X1 i_0_0_533 (.ZN (n_0_0_410), .A (drc_ipo_n33), .B1 (n_0_0_409), .B2 (n_0_0_142));
INV_X1 i_0_0_532 (.ZN (n_0_0_409), .A (n_0_0_321));
NAND2_X1 i_0_0_531 (.ZN (n_0_0_408), .A1 (n_0_0_379), .A2 (drc_ipo_n34));
OAI22_X1 i_0_0_530 (.ZN (n_0_158), .A1 (n_0_0_403), .A2 (n_0_0_109), .B1 (n_0_0_407), .B2 (n_0_0_108));
AOI22_X1 i_0_0_529 (.ZN (n_0_0_407), .A1 (n_0_0_399), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_406));
OAI22_X1 i_0_0_528 (.ZN (n_0_0_406), .A1 (n_0_0_392), .A2 (n_0_0_404), .B1 (n_0_0_292), .B2 (n_0_0_405));
INV_X1 i_0_0_527 (.ZN (n_0_0_405), .A (n_0_0_404));
NOR2_X1 i_0_0_526 (.ZN (n_0_0_404), .A1 (n_0_0_361), .A2 (drc_ipo_n33));
OAI22_X1 i_0_0_525 (.ZN (n_0_157), .A1 (n_0_0_403), .A2 (n_0_0_108), .B1 (n_0_0_400), .B2 (n_0_0_109));
OAI22_X1 i_0_0_524 (.ZN (n_0_0_403), .A1 (n_0_0_396), .A2 (n_0_0_101), .B1 (n_0_0_402), .B2 (hfn_ipo_n32));
OAI21_X1 i_0_0_523 (.ZN (n_0_0_402), .A (n_0_0_401), .B1 (n_0_0_388), .B2 (n_0_0_70));
OAI211_X1 i_0_0_522 (.ZN (n_0_0_401), .A (n_0_0_391), .B (n_0_0_70), .C1 (n_0_0_282), .C2 (n_0_0_361));
OAI22_X1 i_0_0_521 (.ZN (n_0_156), .A1 (n_0_0_397), .A2 (n_0_0_109), .B1 (n_0_0_400), .B2 (n_0_0_108));
AOI22_X1 i_0_0_520 (.ZN (n_0_0_400), .A1 (n_0_0_399), .A2 (n_0_0_101), .B1 (hfn_ipo_n32), .B2 (n_0_0_393));
AOI22_X1 i_0_0_519 (.ZN (n_0_0_399), .A1 (n_0_0_384), .A2 (drc_ipo_n33), .B1 (n_0_0_70), .B2 (n_0_0_398));
OAI21_X1 i_0_0_518 (.ZN (n_0_0_398), .A (n_0_0_391), .B1 (n_0_0_274), .B2 (n_0_0_361));
OAI22_X1 i_0_0_517 (.ZN (n_0_155), .A1 (n_0_0_397), .A2 (n_0_0_108), .B1 (n_0_0_394), .B2 (n_0_0_109));
AOI22_X1 i_0_0_516 (.ZN (n_0_0_397), .A1 (n_0_0_389), .A2 (hfn_ipo_n32), .B1 (n_0_0_396), .B2 (n_0_0_101));
AOI22_X1 i_0_0_515 (.ZN (n_0_0_396), .A1 (n_0_0_380), .A2 (drc_ipo_n33), .B1 (n_0_0_395), .B2 (n_0_0_70));
OAI21_X1 i_0_0_514 (.ZN (n_0_0_395), .A (n_0_0_391), .B1 (n_0_0_265), .B2 (n_0_0_361));
OAI22_X1 i_0_0_513 (.ZN (n_0_154), .A1 (n_0_0_390), .A2 (n_0_0_109), .B1 (n_0_0_394), .B2 (n_0_0_108));
AOI22_X1 i_0_0_512 (.ZN (n_0_0_394), .A1 (n_0_0_385), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_393));
OAI22_X1 i_0_0_511 (.ZN (n_0_0_393), .A1 (n_0_0_376), .A2 (n_0_0_70), .B1 (n_0_0_392), .B2 (drc_ipo_n33));
OAI21_X1 i_0_0_510 (.ZN (n_0_0_392), .A (n_0_0_391), .B1 (n_0_0_255), .B2 (n_0_0_361));
NAND2_X1 i_0_0_509 (.ZN (n_0_0_391), .A1 (n_0_0_321), .A2 (n_0_0_361));
OAI22_X1 i_0_0_508 (.ZN (n_0_153), .A1 (n_0_0_390), .A2 (n_0_0_108), .B1 (n_0_0_386), .B2 (n_0_0_109));
AOI22_X1 i_0_0_507 (.ZN (n_0_0_390), .A1 (hfn_ipo_n32), .A2 (n_0_0_381), .B1 (n_0_0_389), .B2 (n_0_0_101));
OAI22_X1 i_0_0_506 (.ZN (n_0_0_389), .A1 (n_0_0_372), .A2 (n_0_0_70), .B1 (n_0_0_388), .B2 (drc_ipo_n33));
OAI22_X1 i_0_0_505 (.ZN (n_0_0_388), .A1 (n_0_0_356), .A2 (n_0_0_142), .B1 (n_0_0_331), .B2 (n_0_0_387));
NOR2_X1 i_0_0_504 (.ZN (n_0_0_387), .A1 (n_0_0_315), .A2 (n_0_0_69));
OAI22_X1 i_0_0_503 (.ZN (n_0_152), .A1 (n_0_0_382), .A2 (n_0_0_109), .B1 (n_0_0_386), .B2 (n_0_0_108));
AOI22_X1 i_0_0_502 (.ZN (n_0_0_386), .A1 (n_0_0_385), .A2 (n_0_0_101), .B1 (hfn_ipo_n32), .B2 (n_0_0_377));
OAI22_X1 i_0_0_501 (.ZN (n_0_0_385), .A1 (n_0_0_384), .A2 (drc_ipo_n33), .B1 (n_0_0_369), .B2 (n_0_0_70));
OAI22_X1 i_0_0_500 (.ZN (n_0_0_384), .A1 (n_0_0_352), .A2 (n_0_0_142), .B1 (n_0_0_383), .B2 (drc_ipo_n34));
OAI21_X1 i_0_0_499 (.ZN (n_0_0_383), .A (n_0_0_323), .B1 (n_0_0_69), .B2 (n_0_0_307));
OAI22_X1 i_0_0_498 (.ZN (n_0_151), .A1 (n_0_0_382), .A2 (n_0_0_108), .B1 (n_0_0_378), .B2 (n_0_0_109));
OAI22_X1 i_0_0_497 (.ZN (n_0_0_382), .A1 (n_0_0_381), .A2 (hfn_ipo_n32), .B1 (n_0_0_373), .B2 (n_0_0_101));
OAI22_X1 i_0_0_496 (.ZN (n_0_0_381), .A1 (drc_ipo_n33), .A2 (n_0_0_380), .B1 (n_0_0_366), .B2 (n_0_0_70));
OAI22_X1 i_0_0_495 (.ZN (n_0_0_380), .A1 (n_0_0_348), .A2 (n_0_0_142), .B1 (n_0_0_379), .B2 (drc_ipo_n34));
OAI21_X1 i_0_0_494 (.ZN (n_0_0_379), .A (n_0_0_323), .B1 (n_0_0_69), .B2 (n_0_0_299));
OAI22_X1 i_0_0_493 (.ZN (n_0_150), .A1 (n_0_0_374), .A2 (n_0_0_109), .B1 (n_0_0_378), .B2 (n_0_0_108));
OAI22_X1 i_0_0_492 (.ZN (n_0_0_378), .A1 (n_0_0_370), .A2 (n_0_0_101), .B1 (n_0_0_377), .B2 (hfn_ipo_n32));
OAI22_X1 i_0_0_491 (.ZN (n_0_0_377), .A1 (n_0_0_363), .A2 (n_0_0_70), .B1 (drc_ipo_n33), .B2 (n_0_0_376));
NOR2_X1 i_0_0_490 (.ZN (n_0_0_376), .A1 (n_0_0_322), .A2 (n_0_0_375));
OAI22_X1 i_0_0_489 (.ZN (n_0_0_375), .A1 (n_0_0_292), .A2 (n_0_0_326), .B1 (n_0_0_227), .B2 (n_0_0_361));
OAI22_X1 i_0_0_488 (.ZN (n_0_149), .A1 (n_0_0_371), .A2 (n_0_0_109), .B1 (n_0_0_374), .B2 (n_0_0_108));
OAI22_X1 i_0_0_487 (.ZN (n_0_0_374), .A1 (n_0_0_373), .A2 (hfn_ipo_n32), .B1 (n_0_0_367), .B2 (n_0_0_101));
AOI22_X1 i_0_0_486 (.ZN (n_0_0_373), .A1 (n_0_0_372), .A2 (n_0_0_70), .B1 (n_0_0_357), .B2 (drc_ipo_n33));
AOI221_X1 i_0_0_485 (.ZN (n_0_0_372), .A (n_0_0_322), .B1 (n_0_0_218), .B2 (n_0_0_362)
    , .C1 (n_0_0_282), .C2 (n_0_0_344));
OAI22_X1 i_0_0_484 (.ZN (n_0_148), .A1 (n_0_0_371), .A2 (n_0_0_108), .B1 (n_0_0_368), .B2 (n_0_0_109));
OAI22_X1 i_0_0_483 (.ZN (n_0_0_371), .A1 (n_0_0_364), .A2 (n_0_0_101), .B1 (hfn_ipo_n32), .B2 (n_0_0_370));
AOI22_X1 i_0_0_482 (.ZN (n_0_0_370), .A1 (n_0_0_369), .A2 (n_0_0_70), .B1 (n_0_0_353), .B2 (drc_ipo_n33));
AOI221_X1 i_0_0_481 (.ZN (n_0_0_369), .A (n_0_0_322), .B1 (n_0_0_210), .B2 (n_0_0_362)
    , .C1 (n_0_0_274), .C2 (n_0_0_344));
OAI22_X1 i_0_0_480 (.ZN (n_0_147), .A1 (n_0_0_365), .A2 (n_0_0_109), .B1 (n_0_0_368), .B2 (n_0_0_108));
OAI22_X1 i_0_0_479 (.ZN (n_0_0_368), .A1 (n_0_0_367), .A2 (hfn_ipo_n32), .B1 (n_0_0_358), .B2 (n_0_0_101));
AOI22_X1 i_0_0_478 (.ZN (n_0_0_367), .A1 (n_0_0_366), .A2 (n_0_0_70), .B1 (n_0_0_349), .B2 (drc_ipo_n33));
AOI221_X1 i_0_0_477 (.ZN (n_0_0_366), .A (n_0_0_322), .B1 (n_0_0_199), .B2 (n_0_0_362)
    , .C1 (n_0_0_265), .C2 (n_0_0_344));
OAI22_X1 i_0_0_476 (.ZN (n_0_146), .A1 (n_0_0_365), .A2 (n_0_0_108), .B1 (n_0_0_359), .B2 (n_0_0_109));
OAI22_X1 i_0_0_475 (.ZN (n_0_0_365), .A1 (n_0_0_364), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_354));
OAI22_X1 i_0_0_474 (.ZN (n_0_0_364), .A1 (n_0_0_345), .A2 (n_0_0_70), .B1 (drc_ipo_n33), .B2 (n_0_0_363));
AOI21_X1 i_0_0_473 (.ZN (n_0_0_363), .A (n_0_0_360), .B1 (n_0_0_191), .B2 (n_0_0_362));
INV_X1 i_0_0_472 (.ZN (n_0_0_362), .A (n_0_0_361));
NAND2_X1 i_0_0_471 (.ZN (n_0_0_361), .A1 (\shift[4] ), .A2 (drc_ipo_n34));
OAI21_X1 i_0_0_470 (.ZN (n_0_0_360), .A (n_0_0_323), .B1 (n_0_0_256), .B2 (n_0_0_326));
OAI22_X1 i_0_0_469 (.ZN (n_0_145), .A1 (n_0_0_355), .A2 (n_0_0_109), .B1 (n_0_0_359), .B2 (n_0_0_108));
OAI22_X1 i_0_0_468 (.ZN (n_0_0_359), .A1 (n_0_0_350), .A2 (n_0_0_101), .B1 (n_0_0_358), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_0_467 (.ZN (n_0_0_358), .A1 (n_0_0_357), .A2 (n_0_0_70), .B1 (n_0_0_341), .B2 (drc_ipo_n33));
OAI22_X1 i_0_0_466 (.ZN (n_0_0_357), .A1 (n_0_0_356), .A2 (drc_ipo_n34), .B1 (n_0_0_317), .B2 (n_0_0_142));
OAI21_X1 i_0_0_465 (.ZN (n_0_0_356), .A (n_0_0_323), .B1 (n_0_0_69), .B2 (n_0_0_248));
OAI22_X1 i_0_0_464 (.ZN (n_0_144), .A1 (n_0_0_355), .A2 (n_0_0_108), .B1 (n_0_0_351), .B2 (n_0_0_109));
AOI22_X1 i_0_0_463 (.ZN (n_0_0_355), .A1 (n_0_0_346), .A2 (hfn_ipo_n32), .B1 (n_0_0_101), .B2 (n_0_0_354));
AOI22_X1 i_0_0_462 (.ZN (n_0_0_354), .A1 (n_0_0_353), .A2 (n_0_0_70), .B1 (n_0_0_337), .B2 (drc_ipo_n33));
OAI22_X1 i_0_0_461 (.ZN (n_0_0_353), .A1 (n_0_0_352), .A2 (drc_ipo_n34), .B1 (n_0_0_142), .B2 (n_0_0_309));
OAI21_X1 i_0_0_460 (.ZN (n_0_0_352), .A (n_0_0_323), .B1 (n_0_0_69), .B2 (n_0_0_241));
OAI22_X1 i_0_0_459 (.ZN (n_0_143), .A1 (n_0_0_347), .A2 (n_0_0_109), .B1 (n_0_0_351), .B2 (n_0_0_108));
AOI22_X1 i_0_0_458 (.ZN (n_0_0_351), .A1 (n_0_0_350), .A2 (n_0_0_101), .B1 (n_0_0_342), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_0_457 (.ZN (n_0_0_350), .A1 (n_0_0_349), .A2 (n_0_0_70), .B1 (n_0_0_333), .B2 (drc_ipo_n33));
OAI22_X1 i_0_0_456 (.ZN (n_0_0_349), .A1 (n_0_0_348), .A2 (drc_ipo_n34), .B1 (n_0_0_142), .B2 (n_0_0_301));
OAI21_X1 i_0_0_455 (.ZN (n_0_0_348), .A (n_0_0_323), .B1 (n_0_0_69), .B2 (n_0_0_234));
OAI22_X1 i_0_0_454 (.ZN (n_0_142), .A1 (n_0_0_347), .A2 (n_0_0_108), .B1 (n_0_0_343), .B2 (n_0_0_109));
AOI22_X1 i_0_0_453 (.ZN (n_0_0_347), .A1 (n_0_0_346), .A2 (n_0_0_101), .B1 (hfn_ipo_n32), .B2 (n_0_0_338));
OAI22_X1 i_0_0_452 (.ZN (n_0_0_346), .A1 (n_0_0_345), .A2 (drc_ipo_n33), .B1 (n_0_0_328), .B2 (n_0_0_70));
AOI221_X1 i_0_0_451 (.ZN (n_0_0_345), .A (n_0_0_324), .B1 (n_0_0_226), .B2 (n_0_0_344)
    , .C1 (drc_ipo_n34), .C2 (n_0_0_293));
INV_X1 i_0_0_450 (.ZN (n_0_0_344), .A (n_0_0_326));
OAI22_X1 i_0_0_449 (.ZN (n_0_141), .A1 (n_0_0_339), .A2 (n_0_0_109), .B1 (n_0_0_343), .B2 (n_0_0_108));
AOI22_X1 i_0_0_448 (.ZN (n_0_0_343), .A1 (n_0_0_101), .A2 (n_0_0_342), .B1 (n_0_0_334), .B2 (hfn_ipo_n32));
OAI22_X1 i_0_0_447 (.ZN (n_0_0_342), .A1 (n_0_0_341), .A2 (drc_ipo_n33), .B1 (n_0_0_318), .B2 (n_0_0_70));
OAI22_X1 i_0_0_446 (.ZN (n_0_0_341), .A1 (n_0_0_331), .A2 (n_0_0_340), .B1 (n_0_0_142), .B2 (n_0_0_285));
NOR2_X1 i_0_0_445 (.ZN (n_0_0_340), .A1 (n_0_0_219), .A2 (n_0_0_69));
OAI22_X1 i_0_0_444 (.ZN (n_0_140), .A1 (n_0_0_339), .A2 (n_0_0_108), .B1 (n_0_0_335), .B2 (n_0_0_109));
AOI22_X1 i_0_0_443 (.ZN (n_0_0_339), .A1 (n_0_0_329), .A2 (hfn_ipo_n31), .B1 (n_0_0_101), .B2 (n_0_0_338));
OAI22_X1 i_0_0_442 (.ZN (n_0_0_338), .A1 (n_0_0_337), .A2 (drc_ipo_n33), .B1 (n_0_0_310), .B2 (n_0_0_70));
OAI22_X1 i_0_0_441 (.ZN (n_0_0_337), .A1 (n_0_0_331), .A2 (n_0_0_336), .B1 (n_0_0_142), .B2 (n_0_0_276));
NOR2_X1 i_0_0_440 (.ZN (n_0_0_336), .A1 (n_0_0_211), .A2 (n_0_0_69));
OAI22_X1 i_0_0_439 (.ZN (n_0_139), .A1 (n_0_0_330), .A2 (hfn_ipo_n29), .B1 (n_0_0_335), .B2 (n_0_0_108));
AOI22_X1 i_0_0_438 (.ZN (n_0_0_335), .A1 (n_0_0_334), .A2 (n_0_0_101), .B1 (n_0_0_319), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_437 (.ZN (n_0_0_334), .A1 (n_0_0_333), .A2 (drc_ipo_n33), .B1 (n_0_0_70), .B2 (n_0_0_302));
OAI22_X1 i_0_0_436 (.ZN (n_0_0_333), .A1 (n_0_0_331), .A2 (n_0_0_332), .B1 (n_0_0_142), .B2 (n_0_0_267));
NOR2_X1 i_0_0_435 (.ZN (n_0_0_332), .A1 (n_0_0_200), .A2 (n_0_0_69));
NAND2_X1 i_0_0_434 (.ZN (n_0_0_331), .A1 (n_0_0_323), .A2 (n_0_0_142));
OAI22_X1 i_0_0_433 (.ZN (n_0_138), .A1 (n_0_0_330), .A2 (hfn_ipo_n27), .B1 (n_0_0_320), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_432 (.ZN (n_0_0_330), .A1 (n_0_0_329), .A2 (n_0_0_101), .B1 (hfn_ipo_n31), .B2 (n_0_0_311));
OAI22_X1 i_0_0_431 (.ZN (n_0_0_329), .A1 (n_0_0_328), .A2 (drc_ipo_n33), .B1 (n_0_0_294), .B2 (n_0_0_70));
AOI21_X1 i_0_0_430 (.ZN (n_0_0_328), .A (n_0_0_327), .B1 (drc_ipo_n34), .B2 (n_0_0_258));
OAI21_X1 i_0_0_429 (.ZN (n_0_0_327), .A (n_0_0_325), .B1 (n_0_0_192), .B2 (n_0_0_326));
NAND2_X1 i_0_0_428 (.ZN (n_0_0_326), .A1 (n_0_0_142), .A2 (\shift[4] ));
INV_X1 i_0_0_427 (.ZN (n_0_0_325), .A (n_0_0_324));
NOR2_X1 i_0_0_426 (.ZN (n_0_0_324), .A1 (n_0_0_323), .A2 (drc_ipo_n34));
INV_X1 i_0_0_425 (.ZN (n_0_0_323), .A (n_0_0_322));
NOR2_X1 i_0_0_424 (.ZN (n_0_0_322), .A1 (n_0_0_321), .A2 (\shift[4] ));
AOI221_X1 i_0_0_423 (.ZN (n_0_0_321), .A (n_0_0_314), .B1 (n_0_70), .B2 (n_0_0_88)
    , .C1 (\read_data2[31] ), .C2 (n_0_0_89));
OAI22_X1 i_0_0_422 (.ZN (n_0_137), .A1 (n_0_0_320), .A2 (hfn_ipo_n27), .B1 (n_0_0_312), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_421 (.ZN (n_0_0_320), .A1 (n_0_0_319), .A2 (n_0_0_101), .B1 (n_0_0_303), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_420 (.ZN (n_0_0_319), .A1 (n_0_0_318), .A2 (drc_ipo_n33), .B1 (n_0_0_286), .B2 (n_0_0_70));
AOI22_X1 i_0_0_419 (.ZN (n_0_0_318), .A1 (n_0_0_317), .A2 (n_0_0_142), .B1 (drc_ipo_n34), .B2 (n_0_0_249));
OAI22_X1 i_0_0_418 (.ZN (n_0_0_317), .A1 (n_0_0_315), .A2 (\shift[4] ), .B1 (n_0_0_316), .B2 (n_0_0_69));
INV_X1 i_0_0_417 (.ZN (n_0_0_316), .A (n_0_0_185));
AOI221_X1 i_0_0_416 (.ZN (n_0_0_315), .A (n_0_0_314), .B1 (n_0_69), .B2 (n_0_0_88)
    , .C1 (\read_data2[30] ), .C2 (n_0_0_89));
INV_X1 i_0_0_415 (.ZN (n_0_0_314), .A (n_0_0_313));
AOI22_X1 i_0_0_414 (.ZN (n_0_0_313), .A1 (n_0_0_85), .A2 (n_0_39), .B1 (n_0_0_86), .B2 (\read_data2[31] ));
OAI22_X1 i_0_0_413 (.ZN (n_0_136), .A1 (n_0_0_312), .A2 (hfn_ipo_n27), .B1 (n_0_0_304), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_412 (.ZN (n_0_0_312), .A1 (n_0_0_311), .A2 (hfn_ipo_n25), .B1 (n_0_0_295), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_411 (.ZN (n_0_0_311), .A1 (n_0_0_277), .A2 (n_0_0_70), .B1 (n_0_0_310), .B2 (drc_ipo_n33));
AOI22_X1 i_0_0_410 (.ZN (n_0_0_310), .A1 (n_0_0_309), .A2 (n_0_0_142), .B1 (n_0_0_242), .B2 (drc_ipo_n34));
OAI22_X1 i_0_0_409 (.ZN (n_0_0_309), .A1 (n_0_0_307), .A2 (\shift[4] ), .B1 (n_0_0_308), .B2 (n_0_0_69));
INV_X1 i_0_0_408 (.ZN (n_0_0_308), .A (n_0_0_179));
AND2_X1 i_0_0_407 (.ZN (n_0_0_307), .A1 (n_0_0_305), .A2 (n_0_0_306));
AOI22_X1 i_0_0_406 (.ZN (n_0_0_306), .A1 (n_0_0_86), .A2 (\read_data2[30] ), .B1 (\read_data2[29] ), .B2 (n_0_0_89));
AOI22_X1 i_0_0_405 (.ZN (n_0_0_305), .A1 (n_0_0_85), .A2 (n_0_38), .B1 (n_0_0_88), .B2 (n_0_68));
OAI22_X1 i_0_0_404 (.ZN (n_0_135), .A1 (n_0_0_304), .A2 (hfn_ipo_n27), .B1 (n_0_0_296), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_403 (.ZN (n_0_0_304), .A1 (n_0_0_303), .A2 (hfn_ipo_n25), .B1 (n_0_0_287), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_402 (.ZN (n_0_0_303), .A1 (n_0_0_302), .A2 (drc_ipo_n33), .B1 (n_0_0_268), .B2 (n_0_0_70));
AOI22_X1 i_0_0_401 (.ZN (n_0_0_302), .A1 (n_0_0_301), .A2 (n_0_0_142), .B1 (n_0_0_235), .B2 (drc_ipo_n34));
OAI22_X1 i_0_0_400 (.ZN (n_0_0_301), .A1 (n_0_0_299), .A2 (\shift[4] ), .B1 (n_0_0_300), .B2 (n_0_0_69));
INV_X1 i_0_0_399 (.ZN (n_0_0_300), .A (n_0_0_173));
AND2_X1 i_0_0_398 (.ZN (n_0_0_299), .A1 (n_0_0_297), .A2 (n_0_0_298));
AOI22_X1 i_0_0_397 (.ZN (n_0_0_298), .A1 (n_0_0_88), .A2 (n_0_67), .B1 (n_0_0_89), .B2 (\read_data2[28] ));
AOI22_X1 i_0_0_396 (.ZN (n_0_0_297), .A1 (n_0_0_85), .A2 (n_0_37), .B1 (n_0_0_86), .B2 (\read_data2[29] ));
OAI22_X1 i_0_0_395 (.ZN (n_0_134), .A1 (n_0_0_288), .A2 (hfn_ipo_n29), .B1 (n_0_0_296), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_394 (.ZN (n_0_0_296), .A1 (hfn_ipo_n25), .A2 (n_0_0_295), .B1 (n_0_0_278), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_393 (.ZN (n_0_0_295), .A1 (n_0_0_294), .A2 (drc_ipo_n33), .B1 (n_0_0_259), .B2 (n_0_0_70));
AOI22_X1 i_0_0_392 (.ZN (n_0_0_294), .A1 (n_0_0_293), .A2 (n_0_0_142), .B1 (n_0_0_228), .B2 (drc_ipo_n34));
OAI22_X1 i_0_0_391 (.ZN (n_0_0_293), .A1 (n_0_0_289), .A2 (n_0_0_69), .B1 (n_0_0_292), .B2 (\shift[4] ));
AND2_X1 i_0_0_390 (.ZN (n_0_0_292), .A1 (n_0_0_290), .A2 (n_0_0_291));
AOI22_X1 i_0_0_389 (.ZN (n_0_0_291), .A1 (n_0_0_88), .A2 (n_0_66), .B1 (n_0_0_89), .B2 (\read_data2[27] ));
AOI22_X1 i_0_0_388 (.ZN (n_0_0_290), .A1 (n_0_0_85), .A2 (n_0_36), .B1 (n_0_0_86), .B2 (\read_data2[28] ));
INV_X1 i_0_0_387 (.ZN (n_0_0_289), .A (n_0_0_167));
OAI22_X1 i_0_0_386 (.ZN (n_0_133), .A1 (n_0_0_288), .A2 (hfn_ipo_n27), .B1 (n_0_0_279), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_385 (.ZN (n_0_0_288), .A1 (n_0_0_287), .A2 (hfn_ipo_n25), .B1 (n_0_0_269), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_384 (.ZN (n_0_0_287), .A1 (n_0_0_286), .A2 (drc_ipo_n33), .B1 (n_0_0_250), .B2 (n_0_0_70));
AOI22_X1 i_0_0_383 (.ZN (n_0_0_286), .A1 (n_0_0_285), .A2 (n_0_0_142), .B1 (n_0_0_220), .B2 (drc_ipo_n34));
OAI22_X1 i_0_0_382 (.ZN (n_0_0_285), .A1 (n_0_0_283), .A2 (\shift[4] ), .B1 (n_0_0_284), .B2 (n_0_0_69));
INV_X1 i_0_0_381 (.ZN (n_0_0_284), .A (n_0_0_161));
INV_X1 i_0_0_380 (.ZN (n_0_0_283), .A (n_0_0_282));
NAND2_X1 i_0_0_379 (.ZN (n_0_0_282), .A1 (n_0_0_280), .A2 (n_0_0_281));
AOI22_X1 i_0_0_378 (.ZN (n_0_0_281), .A1 (n_0_0_88), .A2 (n_0_65), .B1 (n_0_0_89), .B2 (\read_data2[26] ));
AOI22_X1 i_0_0_377 (.ZN (n_0_0_280), .A1 (n_0_0_85), .A2 (n_0_35), .B1 (n_0_0_86), .B2 (\read_data2[27] ));
OAI22_X1 i_0_0_376 (.ZN (n_0_132), .A1 (n_0_0_279), .A2 (hfn_ipo_n27), .B1 (n_0_0_270), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_375 (.ZN (n_0_0_279), .A1 (n_0_0_278), .A2 (hfn_ipo_n25), .B1 (n_0_0_260), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_374 (.ZN (n_0_0_278), .A1 (n_0_0_277), .A2 (drc_ipo_n33), .B1 (n_0_0_243), .B2 (n_0_0_70));
AOI22_X1 i_0_0_373 (.ZN (n_0_0_277), .A1 (n_0_0_276), .A2 (n_0_0_142), .B1 (n_0_0_212), .B2 (drc_ipo_n34));
OAI22_X1 i_0_0_372 (.ZN (n_0_0_276), .A1 (n_0_0_271), .A2 (n_0_0_69), .B1 (n_0_0_275), .B2 (\shift[4] ));
INV_X1 i_0_0_371 (.ZN (n_0_0_275), .A (n_0_0_274));
NAND2_X1 i_0_0_370 (.ZN (n_0_0_274), .A1 (n_0_0_272), .A2 (n_0_0_273));
AOI22_X1 i_0_0_369 (.ZN (n_0_0_273), .A1 (n_0_0_88), .A2 (n_0_64), .B1 (n_0_0_89), .B2 (\read_data2[25] ));
AOI22_X1 i_0_0_368 (.ZN (n_0_0_272), .A1 (n_0_0_85), .A2 (n_0_34), .B1 (n_0_0_86), .B2 (\read_data2[26] ));
INV_X1 i_0_0_367 (.ZN (n_0_0_271), .A (n_0_0_155));
OAI22_X1 i_0_0_366 (.ZN (n_0_201), .A1 (n_0_0_270), .A2 (hfn_ipo_n27), .B1 (n_0_0_261), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_365 (.ZN (n_0_0_270), .A1 (n_0_0_269), .A2 (hfn_ipo_n25), .B1 (n_0_0_251), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_364 (.ZN (n_0_0_269), .A1 (n_0_0_268), .A2 (drc_ipo_n33), .B1 (n_0_0_236), .B2 (n_0_0_70));
AOI22_X1 i_0_0_363 (.ZN (n_0_0_268), .A1 (n_0_0_201), .A2 (drc_ipo_n34), .B1 (n_0_0_267), .B2 (n_0_0_142));
OAI22_X1 i_0_0_362 (.ZN (n_0_0_267), .A1 (n_0_0_262), .A2 (n_0_0_69), .B1 (n_0_0_266), .B2 (\shift[4] ));
INV_X1 i_0_0_361 (.ZN (n_0_0_266), .A (n_0_0_265));
NAND2_X1 i_0_0_360 (.ZN (n_0_0_265), .A1 (n_0_0_263), .A2 (n_0_0_264));
AOI22_X1 i_0_0_359 (.ZN (n_0_0_264), .A1 (n_0_0_88), .A2 (n_0_63), .B1 (n_0_0_89), .B2 (\read_data2[24] ));
AOI22_X1 i_0_0_358 (.ZN (n_0_0_263), .A1 (n_0_0_85), .A2 (n_0_33), .B1 (n_0_0_86), .B2 (\read_data2[25] ));
INV_X1 i_0_0_357 (.ZN (n_0_0_262), .A (n_0_0_149));
OAI22_X1 i_0_0_356 (.ZN (n_0_200), .A1 (n_0_0_252), .A2 (hfn_ipo_n29), .B1 (n_0_0_261), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_355 (.ZN (n_0_0_261), .A1 (n_0_0_244), .A2 (hfn_ipo_n31), .B1 (n_0_0_260), .B2 (hfn_ipo_n25));
OAI22_X1 i_0_0_354 (.ZN (n_0_0_260), .A1 (n_0_0_259), .A2 (drc_ipo_n33), .B1 (n_0_0_229), .B2 (n_0_0_70));
OAI22_X1 i_0_0_353 (.ZN (n_0_0_259), .A1 (n_0_0_258), .A2 (drc_ipo_n34), .B1 (n_0_0_193), .B2 (n_0_0_142));
OAI22_X1 i_0_0_352 (.ZN (n_0_0_258), .A1 (n_0_0_256), .A2 (\shift[4] ), .B1 (n_0_0_257), .B2 (n_0_0_69));
INV_X1 i_0_0_351 (.ZN (n_0_0_257), .A (n_0_0_140));
INV_X1 i_0_0_350 (.ZN (n_0_0_256), .A (n_0_0_255));
NAND2_X1 i_0_0_349 (.ZN (n_0_0_255), .A1 (n_0_0_253), .A2 (n_0_0_254));
AOI22_X1 i_0_0_348 (.ZN (n_0_0_254), .A1 (n_0_0_88), .A2 (n_0_62), .B1 (n_0_0_89), .B2 (\read_data2[23] ));
AOI22_X1 i_0_0_347 (.ZN (n_0_0_253), .A1 (n_0_0_85), .A2 (n_0_32), .B1 (n_0_0_86), .B2 (\read_data2[24] ));
OAI22_X1 i_0_0_346 (.ZN (n_0_199), .A1 (n_0_0_252), .A2 (hfn_ipo_n27), .B1 (n_0_0_245), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_345 (.ZN (n_0_0_252), .A1 (n_0_0_237), .A2 (hfn_ipo_n31), .B1 (n_0_0_251), .B2 (hfn_ipo_n25));
OAI22_X1 i_0_0_344 (.ZN (n_0_0_251), .A1 (n_0_0_221), .A2 (n_0_0_70), .B1 (n_0_0_250), .B2 (drc_ipo_n33));
AOI22_X1 i_0_0_343 (.ZN (n_0_0_250), .A1 (n_0_0_249), .A2 (n_0_0_142), .B1 (n_0_0_185), .B2 (n_0_0_143));
OAI22_X1 i_0_0_342 (.ZN (n_0_0_249), .A1 (n_0_0_248), .A2 (\shift[4] ), .B1 (n_0_0_134), .B2 (n_0_0_69));
AND2_X1 i_0_0_341 (.ZN (n_0_0_248), .A1 (n_0_0_246), .A2 (n_0_0_247));
AOI22_X1 i_0_0_340 (.ZN (n_0_0_247), .A1 (n_0_0_88), .A2 (n_0_61), .B1 (n_0_0_89), .B2 (\read_data2[22] ));
AOI22_X1 i_0_0_339 (.ZN (n_0_0_246), .A1 (n_0_0_85), .A2 (n_0_31), .B1 (n_0_0_86), .B2 (\read_data2[23] ));
OAI22_X1 i_0_0_338 (.ZN (n_0_198), .A1 (n_0_0_245), .A2 (hfn_ipo_n27), .B1 (n_0_0_238), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_337 (.ZN (n_0_0_245), .A1 (n_0_0_244), .A2 (hfn_ipo_n25), .B1 (n_0_0_230), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_336 (.ZN (n_0_0_244), .A1 (n_0_0_243), .A2 (drc_ipo_n33), .B1 (n_0_0_213), .B2 (n_0_0_70));
AOI22_X1 i_0_0_335 (.ZN (n_0_0_243), .A1 (n_0_0_242), .A2 (n_0_0_142), .B1 (n_0_0_179), .B2 (n_0_0_143));
OAI22_X1 i_0_0_334 (.ZN (n_0_0_242), .A1 (n_0_0_241), .A2 (\shift[4] ), .B1 (n_0_0_128), .B2 (n_0_0_69));
AND2_X1 i_0_0_333 (.ZN (n_0_0_241), .A1 (n_0_0_239), .A2 (n_0_0_240));
AOI22_X1 i_0_0_332 (.ZN (n_0_0_240), .A1 (n_0_0_88), .A2 (n_0_60), .B1 (n_0_0_89), .B2 (\read_data2[21] ));
AOI22_X1 i_0_0_331 (.ZN (n_0_0_239), .A1 (n_0_0_85), .A2 (n_0_30), .B1 (n_0_0_86), .B2 (\read_data2[22] ));
OAI22_X1 i_0_0_330 (.ZN (n_0_197), .A1 (n_0_0_238), .A2 (hfn_ipo_n27), .B1 (n_0_0_231), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_329 (.ZN (n_0_0_238), .A1 (n_0_0_237), .A2 (hfn_ipo_n25), .B1 (n_0_0_222), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_328 (.ZN (n_0_0_237), .A1 (n_0_0_236), .A2 (drc_ipo_n33), .B1 (n_0_0_202), .B2 (n_0_0_70));
AOI22_X1 i_0_0_327 (.ZN (n_0_0_236), .A1 (n_0_0_235), .A2 (n_0_0_142), .B1 (n_0_0_173), .B2 (n_0_0_143));
OAI22_X1 i_0_0_326 (.ZN (n_0_0_235), .A1 (n_0_0_234), .A2 (\shift[4] ), .B1 (n_0_0_121), .B2 (n_0_0_69));
AND2_X1 i_0_0_325 (.ZN (n_0_0_234), .A1 (n_0_0_232), .A2 (n_0_0_233));
AOI22_X1 i_0_0_324 (.ZN (n_0_0_233), .A1 (n_0_0_88), .A2 (n_0_59), .B1 (n_0_0_89), .B2 (\read_data2[20] ));
AOI22_X1 i_0_0_323 (.ZN (n_0_0_232), .A1 (n_0_0_85), .A2 (n_0_29), .B1 (n_0_0_86), .B2 (\read_data2[21] ));
OAI22_X1 i_0_0_322 (.ZN (n_0_196), .A1 (n_0_0_223), .A2 (hfn_ipo_n29), .B1 (n_0_0_231), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_321 (.ZN (n_0_0_231), .A1 (hfn_ipo_n25), .A2 (n_0_0_230), .B1 (n_0_0_214), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_320 (.ZN (n_0_0_230), .A1 (n_0_0_229), .A2 (drc_ipo_n33), .B1 (n_0_0_194), .B2 (n_0_0_70));
AOI22_X1 i_0_0_319 (.ZN (n_0_0_229), .A1 (n_0_0_228), .A2 (n_0_0_142), .B1 (n_0_0_167), .B2 (n_0_0_143));
OAI22_X1 i_0_0_318 (.ZN (n_0_0_228), .A1 (n_0_0_113), .A2 (n_0_0_69), .B1 (n_0_0_227), .B2 (\shift[4] ));
INV_X1 i_0_0_317 (.ZN (n_0_0_227), .A (n_0_0_226));
NAND2_X1 i_0_0_316 (.ZN (n_0_0_226), .A1 (n_0_0_224), .A2 (n_0_0_225));
AOI22_X1 i_0_0_315 (.ZN (n_0_0_225), .A1 (n_0_0_88), .A2 (n_0_58), .B1 (n_0_0_89), .B2 (\read_data2[19] ));
AOI22_X1 i_0_0_314 (.ZN (n_0_0_224), .A1 (n_0_0_85), .A2 (n_0_28), .B1 (n_0_0_86), .B2 (\read_data2[20] ));
OAI22_X1 i_0_0_313 (.ZN (n_0_195), .A1 (n_0_0_223), .A2 (hfn_ipo_n27), .B1 (n_0_0_215), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_312 (.ZN (n_0_0_223), .A1 (n_0_0_222), .A2 (hfn_ipo_n25), .B1 (n_0_0_203), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_311 (.ZN (n_0_0_222), .A1 (n_0_0_221), .A2 (drc_ipo_n33), .B1 (n_0_0_186), .B2 (n_0_0_114));
AOI22_X1 i_0_0_310 (.ZN (n_0_0_221), .A1 (n_0_0_220), .A2 (n_0_0_142), .B1 (n_0_0_161), .B2 (n_0_0_143));
OAI22_X1 i_0_0_309 (.ZN (n_0_0_220), .A1 (n_0_0_135), .A2 (n_0_0_69), .B1 (n_0_0_219), .B2 (\shift[4] ));
INV_X1 i_0_0_308 (.ZN (n_0_0_219), .A (n_0_0_218));
NAND2_X1 i_0_0_307 (.ZN (n_0_0_218), .A1 (n_0_0_216), .A2 (n_0_0_217));
AOI22_X1 i_0_0_306 (.ZN (n_0_0_217), .A1 (n_0_0_88), .A2 (n_0_57), .B1 (n_0_0_89), .B2 (\read_data2[18] ));
AOI22_X1 i_0_0_305 (.ZN (n_0_0_216), .A1 (n_0_0_85), .A2 (n_0_27), .B1 (n_0_0_86), .B2 (\read_data2[19] ));
AOI22_X1 i_0_0_304 (.ZN (n_0_194), .A1 (n_0_0_207), .A2 (hfn_ipo_n27), .B1 (n_0_0_215), .B2 (n_0_0_93));
AOI22_X1 i_0_0_303 (.ZN (n_0_0_215), .A1 (n_0_0_214), .A2 (hfn_ipo_n25), .B1 (n_0_0_195), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_302 (.ZN (n_0_0_214), .A1 (n_0_0_213), .A2 (drc_ipo_n33), .B1 (n_0_0_70), .B2 (n_0_0_180));
AOI22_X1 i_0_0_301 (.ZN (n_0_0_213), .A1 (n_0_0_212), .A2 (n_0_0_142), .B1 (n_0_0_155), .B2 (n_0_0_143));
OAI22_X1 i_0_0_300 (.ZN (n_0_0_212), .A1 (n_0_0_211), .A2 (\shift[4] ), .B1 (n_0_0_124), .B2 (n_0_0_69));
INV_X1 i_0_0_299 (.ZN (n_0_0_211), .A (n_0_0_210));
NAND2_X1 i_0_0_298 (.ZN (n_0_0_210), .A1 (n_0_0_208), .A2 (n_0_0_209));
AOI22_X1 i_0_0_297 (.ZN (n_0_0_209), .A1 (n_0_0_88), .A2 (n_0_56), .B1 (n_0_0_89), .B2 (\read_data2[17] ));
AOI22_X1 i_0_0_296 (.ZN (n_0_0_208), .A1 (n_0_0_85), .A2 (n_0_26), .B1 (n_0_0_86), .B2 (\read_data2[18] ));
AOI22_X1 i_0_0_295 (.ZN (n_0_193), .A1 (n_0_0_207), .A2 (hfn_ipo_n29), .B1 (\shift[0] ), .B2 (n_0_0_196));
NAND2_X1 i_0_0_294 (.ZN (n_0_0_207), .A1 (n_0_0_206), .A2 (n_0_0_68));
AOI22_X1 i_0_0_293 (.ZN (n_0_0_206), .A1 (n_0_0_204), .A2 (hfn_ipo_n25), .B1 (n_0_0_205), .B2 (hfn_ipo_n31));
INV_X1 i_0_0_292 (.ZN (n_0_0_205), .A (n_0_0_187));
INV_X1 i_0_0_291 (.ZN (n_0_0_204), .A (n_0_0_203));
OAI22_X1 i_0_0_290 (.ZN (n_0_0_203), .A1 (n_0_0_202), .A2 (drc_ipo_n33), .B1 (n_0_0_174), .B2 (n_0_0_114));
AOI22_X1 i_0_0_289 (.ZN (n_0_0_202), .A1 (n_0_0_201), .A2 (n_0_0_142), .B1 (n_0_0_149), .B2 (n_0_0_143));
OAI22_X1 i_0_0_288 (.ZN (n_0_0_201), .A1 (n_0_0_200), .A2 (\shift[4] ), .B1 (n_0_0_92), .B2 (n_0_0_69));
INV_X1 i_0_0_287 (.ZN (n_0_0_200), .A (n_0_0_199));
NAND2_X1 i_0_0_286 (.ZN (n_0_0_199), .A1 (n_0_0_197), .A2 (n_0_0_198));
AOI22_X1 i_0_0_285 (.ZN (n_0_0_198), .A1 (n_0_0_88), .A2 (n_0_55), .B1 (n_0_0_89), .B2 (\read_data2[16] ));
AOI22_X1 i_0_0_284 (.ZN (n_0_0_197), .A1 (n_0_0_85), .A2 (n_0_25), .B1 (n_0_0_86), .B2 (\read_data2[17] ));
OAI22_X1 i_0_0_283 (.ZN (n_0_192), .A1 (n_0_0_196), .A2 (hfn_ipo_n27), .B1 (n_0_0_188), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_282 (.ZN (n_0_0_196), .A1 (n_0_0_195), .A2 (hfn_ipo_n25), .B1 (hfn_ipo_n31), .B2 (n_0_0_181));
OAI22_X1 i_0_0_281 (.ZN (n_0_0_195), .A1 (n_0_0_194), .A2 (drc_ipo_n33), .B1 (n_0_0_168), .B2 (n_0_0_114));
AOI22_X1 i_0_0_280 (.ZN (n_0_0_194), .A1 (n_0_0_193), .A2 (n_0_0_142), .B1 (n_0_0_140), .B2 (n_0_0_143));
AOI22_X1 i_0_0_279 (.ZN (n_0_0_193), .A1 (n_0_0_192), .A2 (n_0_0_69), .B1 (n_0_0_67), .B2 (\shift[4] ));
INV_X1 i_0_0_278 (.ZN (n_0_0_192), .A (n_0_0_191));
NAND2_X1 i_0_0_277 (.ZN (n_0_0_191), .A1 (n_0_0_189), .A2 (n_0_0_190));
AOI22_X1 i_0_0_276 (.ZN (n_0_0_190), .A1 (n_0_0_88), .A2 (n_0_54), .B1 (n_0_0_89), .B2 (\read_data2[15] ));
AOI22_X1 i_0_0_275 (.ZN (n_0_0_189), .A1 (n_0_0_85), .A2 (n_0_24), .B1 (n_0_0_86), .B2 (\read_data2[16] ));
OAI22_X1 i_0_0_274 (.ZN (n_0_191), .A1 (n_0_0_188), .A2 (hfn_ipo_n27), .B1 (n_0_0_182), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_273 (.ZN (n_0_0_188), .A1 (n_0_0_175), .A2 (hfn_ipo_n31), .B1 (n_0_0_187), .B2 (hfn_ipo_n25));
OAI22_X1 i_0_0_272 (.ZN (n_0_0_187), .A1 (n_0_0_162), .A2 (n_0_0_114), .B1 (n_0_0_186), .B2 (n_0_0_71));
AOI22_X1 i_0_0_271 (.ZN (n_0_0_186), .A1 (n_0_0_133), .A2 (drc_ipo_n34), .B1 (n_0_0_185), .B2 (n_0_0_142));
NAND2_X1 i_0_0_270 (.ZN (n_0_0_185), .A1 (n_0_0_183), .A2 (n_0_0_184));
AOI22_X1 i_0_0_269 (.ZN (n_0_0_184), .A1 (n_0_0_88), .A2 (n_0_53), .B1 (n_0_0_89), .B2 (\read_data2[14] ));
AOI22_X1 i_0_0_268 (.ZN (n_0_0_183), .A1 (n_0_0_85), .A2 (n_0_23), .B1 (n_0_0_86), .B2 (\read_data2[15] ));
OAI22_X1 i_0_0_267 (.ZN (n_0_190), .A1 (n_0_0_176), .A2 (hfn_ipo_n29), .B1 (n_0_0_182), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_266 (.ZN (n_0_0_182), .A1 (n_0_0_181), .A2 (hfn_ipo_n25), .B1 (n_0_0_169), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_265 (.ZN (n_0_0_181), .A1 (n_0_0_156), .A2 (n_0_0_114), .B1 (n_0_0_180), .B2 (drc_ipo_n33));
AOI22_X1 i_0_0_264 (.ZN (n_0_0_180), .A1 (n_0_0_179), .A2 (n_0_0_141), .B1 (n_0_0_127), .B2 (n_0_0_143));
NAND2_X1 i_0_0_263 (.ZN (n_0_0_179), .A1 (n_0_0_177), .A2 (n_0_0_178));
AOI22_X1 i_0_0_262 (.ZN (n_0_0_178), .A1 (n_0_0_88), .A2 (n_0_52), .B1 (n_0_0_89), .B2 (\read_data2[13] ));
AOI22_X1 i_0_0_261 (.ZN (n_0_0_177), .A1 (n_0_0_85), .A2 (n_0_22), .B1 (n_0_0_86), .B2 (\read_data2[14] ));
OAI22_X1 i_0_0_260 (.ZN (n_0_189), .A1 (n_0_0_176), .A2 (hfn_ipo_n27), .B1 (n_0_0_170), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_259 (.ZN (n_0_0_176), .A1 (n_0_0_175), .A2 (hfn_ipo_n25), .B1 (n_0_0_163), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_258 (.ZN (n_0_0_175), .A1 (n_0_0_150), .A2 (n_0_0_70), .B1 (n_0_0_174), .B2 (n_0_0_71));
AOI22_X1 i_0_0_257 (.ZN (n_0_0_174), .A1 (n_0_0_120), .A2 (drc_ipo_n34), .B1 (n_0_0_173), .B2 (n_0_0_142));
NAND2_X1 i_0_0_256 (.ZN (n_0_0_173), .A1 (n_0_0_171), .A2 (n_0_0_172));
AOI22_X1 i_0_0_255 (.ZN (n_0_0_172), .A1 (n_0_0_88), .A2 (n_0_51), .B1 (n_0_0_89), .B2 (\read_data2[12] ));
AOI22_X1 i_0_0_254 (.ZN (n_0_0_171), .A1 (n_0_0_85), .A2 (n_0_21), .B1 (n_0_0_86), .B2 (\read_data2[13] ));
OAI22_X1 i_0_0_253 (.ZN (n_0_188), .A1 (n_0_0_164), .A2 (hfn_ipo_n29), .B1 (n_0_0_170), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_252 (.ZN (n_0_0_170), .A1 (hfn_ipo_n25), .A2 (n_0_0_169), .B1 (n_0_0_157), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_251 (.ZN (n_0_0_169), .A1 (n_0_0_168), .A2 (n_0_0_71), .B1 (n_0_0_144), .B2 (n_0_0_70));
AOI22_X1 i_0_0_250 (.ZN (n_0_0_168), .A1 (n_0_0_167), .A2 (n_0_0_142), .B1 (n_0_0_112), .B2 (drc_ipo_n34));
NAND2_X1 i_0_0_249 (.ZN (n_0_0_167), .A1 (n_0_0_165), .A2 (n_0_0_166));
AOI22_X1 i_0_0_248 (.ZN (n_0_0_166), .A1 (n_0_0_88), .A2 (n_0_50), .B1 (n_0_0_89), .B2 (\read_data2[11] ));
AOI22_X1 i_0_0_247 (.ZN (n_0_0_165), .A1 (n_0_0_85), .A2 (n_0_20), .B1 (n_0_0_86), .B2 (\read_data2[12] ));
OAI22_X1 i_0_0_246 (.ZN (n_0_187), .A1 (n_0_0_164), .A2 (hfn_ipo_n27), .B1 (n_0_0_158), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_245 (.ZN (n_0_0_164), .A1 (n_0_0_163), .A2 (hfn_ipo_n25), .B1 (n_0_0_151), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_244 (.ZN (n_0_0_163), .A1 (n_0_0_162), .A2 (n_0_0_71), .B1 (n_0_0_134), .B2 (n_0_0_115));
AOI22_X1 i_0_0_243 (.ZN (n_0_0_162), .A1 (n_0_0_161), .A2 (n_0_0_142), .B1 (n_0_0_106), .B2 (drc_ipo_n34));
NAND2_X1 i_0_0_242 (.ZN (n_0_0_161), .A1 (n_0_0_159), .A2 (n_0_0_160));
AOI22_X1 i_0_0_241 (.ZN (n_0_0_160), .A1 (n_0_0_88), .A2 (n_0_49), .B1 (n_0_0_89), .B2 (\read_data2[10] ));
AOI22_X1 i_0_0_240 (.ZN (n_0_0_159), .A1 (n_0_0_85), .A2 (n_0_19), .B1 (n_0_0_86), .B2 (\read_data2[11] ));
OAI22_X1 i_0_0_239 (.ZN (n_0_186), .A1 (n_0_0_152), .A2 (hfn_ipo_n29), .B1 (n_0_0_158), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_0_238 (.ZN (n_0_0_158), .A1 (n_0_0_157), .A2 (hfn_ipo_n25), .B1 (n_0_0_145), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_237 (.ZN (n_0_0_157), .A1 (n_0_0_156), .A2 (n_0_0_71), .B1 (n_0_0_128), .B2 (n_0_0_115));
AOI22_X1 i_0_0_236 (.ZN (n_0_0_156), .A1 (n_0_0_99), .A2 (drc_ipo_n34), .B1 (n_0_0_155), .B2 (n_0_0_142));
NAND2_X1 i_0_0_235 (.ZN (n_0_0_155), .A1 (n_0_0_153), .A2 (n_0_0_154));
AOI22_X1 i_0_0_234 (.ZN (n_0_0_154), .A1 (n_0_0_88), .A2 (n_0_48), .B1 (n_0_0_89), .B2 (\read_data2[9] ));
AOI22_X1 i_0_0_233 (.ZN (n_0_0_153), .A1 (n_0_0_85), .A2 (n_0_18), .B1 (n_0_0_86), .B2 (\read_data2[10] ));
OAI22_X1 i_0_0_232 (.ZN (n_0_185), .A1 (n_0_0_152), .A2 (hfn_ipo_n27), .B1 (n_0_0_146), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_231 (.ZN (n_0_0_152), .A1 (n_0_0_151), .A2 (hfn_ipo_n25), .B1 (n_0_0_136), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_230 (.ZN (n_0_0_151), .A1 (n_0_0_150), .A2 (drc_ipo_n33), .B1 (n_0_0_121), .B2 (n_0_0_115));
AOI22_X1 i_0_0_229 (.ZN (n_0_0_150), .A1 (n_0_0_91), .A2 (n_0_0_143), .B1 (n_0_0_149), .B2 (n_0_0_141));
NAND2_X1 i_0_0_228 (.ZN (n_0_0_149), .A1 (n_0_0_147), .A2 (n_0_0_148));
AOI22_X1 i_0_0_227 (.ZN (n_0_0_148), .A1 (n_0_0_88), .A2 (n_0_47), .B1 (n_0_0_89), .B2 (\read_data2[8] ));
AOI22_X1 i_0_0_226 (.ZN (n_0_0_147), .A1 (n_0_0_85), .A2 (n_0_17), .B1 (n_0_0_86), .B2 (\read_data2[9] ));
OAI22_X1 i_0_0_225 (.ZN (n_0_184), .A1 (n_0_0_146), .A2 (hfn_ipo_n27), .B1 (n_0_0_137), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_224 (.ZN (n_0_0_146), .A1 (n_0_0_145), .A2 (hfn_ipo_n25), .B1 (n_0_0_129), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_223 (.ZN (n_0_0_145), .A1 (n_0_0_144), .A2 (drc_ipo_n33), .B1 (n_0_0_113), .B2 (n_0_0_115));
AOI22_X1 i_0_0_222 (.ZN (n_0_0_144), .A1 (n_0_0_140), .A2 (n_0_0_141), .B1 (n_0_0_100), .B2 (n_0_0_143));
NOR2_X1 i_0_0_221 (.ZN (n_0_0_143), .A1 (n_0_0_142), .A2 (\shift[4] ));
INV_X4 i_0_0_220 (.ZN (n_0_0_142), .A (drc_ipo_n34));
NOR2_X1 i_0_0_219 (.ZN (n_0_0_141), .A1 (\shift[4] ), .A2 (drc_ipo_n34));
NAND2_X1 i_0_0_218 (.ZN (n_0_0_140), .A1 (n_0_0_138), .A2 (n_0_0_139));
AOI22_X1 i_0_0_217 (.ZN (n_0_0_139), .A1 (n_0_0_88), .A2 (n_0_46), .B1 (n_0_0_89), .B2 (\read_data2[7] ));
AOI22_X1 i_0_0_216 (.ZN (n_0_0_138), .A1 (n_0_0_85), .A2 (n_0_16), .B1 (n_0_0_86), .B2 (\read_data2[8] ));
OAI22_X1 i_0_0_215 (.ZN (n_0_183), .A1 (n_0_0_137), .A2 (hfn_ipo_n27), .B1 (n_0_0_130), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_214 (.ZN (n_0_0_137), .A1 (n_0_0_122), .A2 (hfn_ipo_n31), .B1 (n_0_0_136), .B2 (hfn_ipo_n25));
OAI22_X1 i_0_0_213 (.ZN (n_0_0_136), .A1 (n_0_0_134), .A2 (n_0_0_72), .B1 (n_0_0_135), .B2 (n_0_0_115));
INV_X1 i_0_0_212 (.ZN (n_0_0_135), .A (n_0_0_106));
INV_X1 i_0_0_211 (.ZN (n_0_0_134), .A (n_0_0_133));
NAND2_X1 i_0_0_210 (.ZN (n_0_0_133), .A1 (n_0_0_131), .A2 (n_0_0_132));
AOI22_X1 i_0_0_209 (.ZN (n_0_0_132), .A1 (n_0_0_88), .A2 (n_0_45), .B1 (n_0_0_89), .B2 (\read_data2[6] ));
AOI22_X1 i_0_0_208 (.ZN (n_0_0_131), .A1 (n_0_0_85), .A2 (n_0_15), .B1 (n_0_0_86), .B2 (\read_data2[7] ));
OAI22_X1 i_0_0_207 (.ZN (n_0_182), .A1 (n_0_0_130), .A2 (hfn_ipo_n27), .B1 (n_0_0_123), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_206 (.ZN (n_0_0_130), .A1 (n_0_0_129), .A2 (hfn_ipo_n25), .B1 (n_0_0_116), .B2 (hfn_ipo_n31));
OAI22_X1 i_0_0_205 (.ZN (n_0_0_129), .A1 (n_0_0_124), .A2 (n_0_0_115), .B1 (n_0_0_128), .B2 (n_0_0_72));
INV_X1 i_0_0_204 (.ZN (n_0_0_128), .A (n_0_0_127));
NAND2_X1 i_0_0_203 (.ZN (n_0_0_127), .A1 (n_0_0_125), .A2 (n_0_0_126));
AOI22_X1 i_0_0_202 (.ZN (n_0_0_126), .A1 (n_0_0_88), .A2 (n_0_44), .B1 (n_0_0_89), .B2 (\read_data2[5] ));
AOI22_X1 i_0_0_201 (.ZN (n_0_0_125), .A1 (n_0_0_85), .A2 (n_0_14), .B1 (n_0_0_86), .B2 (\read_data2[6] ));
INV_X1 i_0_0_200 (.ZN (n_0_0_124), .A (n_0_0_99));
OAI22_X1 i_0_0_199 (.ZN (n_0_181), .A1 (n_0_0_123), .A2 (hfn_ipo_n27), .B1 (n_0_0_117), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_0_198 (.ZN (n_0_0_123), .A1 (n_0_0_122), .A2 (hfn_ipo_n25), .B1 (n_0_0_106), .B2 (n_0_0_102));
OAI22_X1 i_0_0_197 (.ZN (n_0_0_122), .A1 (n_0_0_121), .A2 (n_0_0_72), .B1 (n_0_0_92), .B2 (n_0_0_115));
INV_X1 i_0_0_196 (.ZN (n_0_0_121), .A (n_0_0_120));
NAND2_X1 i_0_0_195 (.ZN (n_0_0_120), .A1 (n_0_0_118), .A2 (n_0_0_119));
AOI22_X1 i_0_0_194 (.ZN (n_0_0_119), .A1 (n_0_0_88), .A2 (n_0_43), .B1 (n_0_0_89), .B2 (\read_data2[4] ));
AOI22_X1 i_0_0_193 (.ZN (n_0_0_118), .A1 (n_0_0_85), .A2 (n_0_13), .B1 (n_0_0_86), .B2 (\read_data2[5] ));
OAI22_X1 i_0_0_192 (.ZN (n_0_180), .A1 (n_0_0_117), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n29), .B2 (n_0_0_107));
AOI22_X1 i_0_0_191 (.ZN (n_0_0_117), .A1 (n_0_0_116), .A2 (hfn_ipo_n25), .B1 (n_0_0_99), .B2 (n_0_0_102));
OAI22_X1 i_0_0_190 (.ZN (n_0_0_116), .A1 (n_0_0_113), .A2 (n_0_0_72), .B1 (n_0_0_67), .B2 (n_0_0_115));
OR2_X1 i_0_0_189 (.ZN (n_0_0_115), .A1 (n_0_0_114), .A2 (drc_ipo_n34));
NAND2_X1 i_0_0_188 (.ZN (n_0_0_114), .A1 (n_0_0_69), .A2 (drc_ipo_n33));
INV_X1 i_0_0_187 (.ZN (n_0_0_113), .A (n_0_0_112));
NAND2_X1 i_0_0_186 (.ZN (n_0_0_112), .A1 (n_0_0_110), .A2 (n_0_0_111));
AOI22_X1 i_0_0_185 (.ZN (n_0_0_111), .A1 (n_0_0_88), .A2 (n_0_42), .B1 (n_0_0_89), .B2 (\read_data2[3] ));
AOI22_X1 i_0_0_184 (.ZN (n_0_0_110), .A1 (n_0_0_85), .A2 (n_0_12), .B1 (n_0_0_86), .B2 (\read_data2[4] ));
OAI22_X1 i_0_0_183 (.ZN (n_0_179), .A1 (n_0_0_107), .A2 (hfn_ipo_n27), .B1 (n_0_0_103), .B2 (hfn_ipo_n29));
NAND2_X1 i_0_0_182 (.ZN (n_0_0_109), .A1 (n_0_0_68), .A2 (\shift[0] ));
INV_X1 i_0_0_181 (.ZN (n_0_0_108), .A (n_0_0_95));
AOI22_X1 i_0_0_180 (.ZN (n_0_0_107), .A1 (n_0_0_91), .A2 (n_0_0_102), .B1 (n_0_0_106), .B2 (n_0_0_73));
NAND2_X1 i_0_0_179 (.ZN (n_0_0_106), .A1 (n_0_0_104), .A2 (n_0_0_105));
AOI22_X1 i_0_0_178 (.ZN (n_0_0_105), .A1 (n_0_0_88), .A2 (n_0_41), .B1 (n_0_0_89), .B2 (\read_data2[2] ));
AOI22_X1 i_0_0_177 (.ZN (n_0_0_104), .A1 (n_0_0_85), .A2 (n_0_11), .B1 (n_0_0_86), .B2 (\read_data2[3] ));
AOI21_X1 i_0_0_176 (.ZN (n_0_178), .A (n_0_0_96), .B1 (n_0_0_103), .B2 (n_0_0_93));
AOI22_X1 i_0_0_175 (.ZN (n_0_0_103), .A1 (n_0_0_99), .A2 (n_0_0_73), .B1 (n_0_0_100), .B2 (n_0_0_102));
NOR2_X1 i_0_0_174 (.ZN (n_0_0_102), .A1 (n_0_0_72), .A2 (hfn_ipo_n25));
INV_X1 i_0_0_173 (.ZN (n_0_0_101), .A (hfn_ipo_n32));
INV_X1 i_0_0_172 (.ZN (n_0_0_100), .A (n_0_0_67));
NAND2_X1 i_0_0_171 (.ZN (n_0_0_99), .A1 (n_0_0_97), .A2 (n_0_0_98));
AOI22_X1 i_0_0_170 (.ZN (n_0_0_98), .A1 (n_0_0_88), .A2 (n_0_40), .B1 (n_0_0_89), .B2 (\read_data2[1] ));
AOI22_X1 i_0_0_169 (.ZN (n_0_0_97), .A1 (n_0_0_85), .A2 (n_0_10), .B1 (n_0_0_86), .B2 (\read_data2[2] ));
AOI21_X1 i_0_0_168 (.ZN (n_0_0_96), .A (n_0_0_95), .B1 (n_0_0_91), .B2 (n_0_0_74));
NOR2_X1 i_0_0_167 (.ZN (n_0_0_95), .A1 (n_0_0_94), .A2 (\shift[0] ));
INV_X1 i_0_0_166 (.ZN (n_0_0_94), .A (n_0_0_68));
AOI221_X1 i_0_0_165 (.ZN (n_0_177), .A (n_0_0_75), .B1 (\shift[0] ), .B2 (n_0_0_67)
    , .C1 (n_0_0_92), .C2 (n_0_0_93));
INV_X1 i_0_0_164 (.ZN (n_0_0_93), .A (\shift[0] ));
INV_X1 i_0_0_163 (.ZN (n_0_0_92), .A (n_0_0_91));
NAND2_X1 i_0_0_162 (.ZN (n_0_0_91), .A1 (n_0_0_87), .A2 (n_0_0_90));
OAI21_X1 i_0_0_161 (.ZN (n_0_0_90), .A (\read_data2[0] ), .B1 (n_0_0_88), .B2 (n_0_0_89));
NOR2_X4 i_0_0_160 (.ZN (n_0_0_89), .A1 (n_0_0_84), .A2 (n_0_0_64));
NOR2_X4 i_0_0_159 (.ZN (n_0_0_88), .A1 (n_0_0_63), .A2 (n_0_0_83));
AOI22_X1 i_0_0_158 (.ZN (n_0_0_87), .A1 (n_0_0_85), .A2 (n_0_9), .B1 (n_0_0_86), .B2 (\read_data2[1] ));
NOR2_X4 i_0_0_157 (.ZN (n_0_0_86), .A1 (n_0_0_65), .A2 (n_0_0_84));
AND3_X2 i_0_0_156 (.ZN (n_0_0_85), .A1 (n_0_0_84), .A2 (n_0_0_64), .A3 (n_0_0_63));
INV_X1 i_0_0_155 (.ZN (n_0_0_84), .A (n_0_0_83));
AOI21_X1 i_0_0_154 (.ZN (n_0_0_83), .A (n_0_0_81), .B1 (n_0_0_16), .B2 (n_0_0_82));
INV_X1 i_0_0_153 (.ZN (n_0_0_82), .A (n_0_0_55));
AOI221_X1 i_0_0_152 (.ZN (n_0_0_81), .A (n_0_0_16), .B1 (n_0_0_79), .B2 (\i[1] ), .C1 (n_0_0_80), .C2 (n_0_0_18));
INV_X1 i_0_0_151 (.ZN (n_0_0_80), .A (n_0_0_38));
AOI21_X1 i_0_0_150 (.ZN (n_0_0_79), .A (n_0_0_78), .B1 (n_0_0_25), .B2 (n_0_0_23));
OAI21_X1 i_0_0_149 (.ZN (n_0_0_78), .A (n_0_0_76), .B1 (n_0_0_25), .B2 (n_0_0_77));
AOI22_X1 i_0_0_148 (.ZN (n_0_0_77), .A1 (n_0_0_19), .A2 (\read_data[31] ), .B1 (n_0_0_20), .B2 (\read_data[23] ));
OAI221_X1 i_0_0_147 (.ZN (n_0_0_76), .A (n_0_0_30), .B1 (\i[3] ), .B2 (\read_data[7] )
    , .C1 (n_0_0_14), .C2 (\read_data[15] ));
NOR3_X1 i_0_0_146 (.ZN (n_0_176), .A1 (n_0_0_67), .A2 (\shift[0] ), .A3 (n_0_0_75));
INV_X1 i_0_0_145 (.ZN (n_0_0_75), .A (n_0_0_74));
AND2_X1 i_0_0_144 (.ZN (n_0_0_74), .A1 (n_0_0_68), .A2 (n_0_0_73));
NOR2_X1 i_0_0_143 (.ZN (n_0_0_73), .A1 (n_0_0_72), .A2 (hfn_ipo_n31));
OR2_X1 i_0_0_142 (.ZN (n_0_0_72), .A1 (n_0_0_71), .A2 (drc_ipo_n34));
NAND2_X1 i_0_0_141 (.ZN (n_0_0_71), .A1 (n_0_0_69), .A2 (n_0_0_70));
INV_X4 i_0_0_140 (.ZN (n_0_0_70), .A (drc_ipo_n33));
INV_X1 i_0_0_139 (.ZN (n_0_0_69), .A (\shift[4] ));
NOR2_X1 i_0_0_138 (.ZN (n_0_0_68), .A1 (n_0_0_17), .A2 (start));
NAND2_X1 i_0_0_137 (.ZN (n_0_0_67), .A1 (n_0_0_66), .A2 (\read_data2[0] ));
INV_X1 i_0_0_136 (.ZN (n_0_0_66), .A (n_0_0_65));
NAND2_X1 i_0_0_135 (.ZN (n_0_0_65), .A1 (n_0_0_63), .A2 (n_0_0_64));
NAND2_X1 i_0_0_134 (.ZN (n_0_0_64), .A1 (n_0_0_56), .A2 (n_0_0_62));
OR2_X1 i_0_0_133 (.ZN (n_0_0_63), .A1 (n_0_0_56), .A2 (n_0_0_62));
AOI22_X1 i_0_0_132 (.ZN (n_0_0_62), .A1 (n_0_0_39), .A2 (\i[0] ), .B1 (n_0_0_61), .B2 (n_0_0_16));
OAI21_X1 i_0_0_131 (.ZN (n_0_0_61), .A (n_0_0_57), .B1 (n_0_0_60), .B2 (\i[1] ));
AOI22_X1 i_0_0_130 (.ZN (n_0_0_60), .A1 (n_0_0_51), .A2 (\i[2] ), .B1 (n_0_0_59), .B2 (n_0_0_25));
AOI221_X1 i_0_0_129 (.ZN (n_0_0_59), .A (n_0_0_58), .B1 (n_0_0_19), .B2 (\read_data[22] )
    , .C1 (\read_data[14] ), .C2 (n_0_0_20));
AND3_X1 i_0_0_128 (.ZN (n_0_0_58), .A1 (n_0_0_26), .A2 (\read_data[6] ), .A3 (\i[3] ));
OR3_X1 i_0_0_127 (.ZN (n_0_0_57), .A1 (n_0_0_44), .A2 (n_0_0_18), .A3 (n_0_0_46));
OAI22_X1 i_0_0_126 (.ZN (n_0_0_56), .A1 (n_0_0_39), .A2 (\i[0] ), .B1 (n_0_0_55), .B2 (n_0_0_16));
OAI21_X1 i_0_0_125 (.ZN (n_0_0_55), .A (n_0_0_47), .B1 (n_0_0_52), .B2 (n_0_0_54));
NAND2_X1 i_0_0_124 (.ZN (n_0_0_54), .A1 (n_0_0_53), .A2 (\i[1] ));
OAI221_X1 i_0_0_123 (.ZN (n_0_0_53), .A (n_0_0_30), .B1 (\read_data[6] ), .B2 (\i[3] )
    , .C1 (n_0_0_14), .C2 (\read_data[14] ));
AOI21_X1 i_0_0_122 (.ZN (n_0_0_52), .A (n_0_0_48), .B1 (n_0_0_51), .B2 (n_0_0_25));
AOI221_X1 i_0_0_121 (.ZN (n_0_0_51), .A (n_0_0_50), .B1 (\read_data[26] ), .B2 (n_0_0_19)
    , .C1 (\read_data[18] ), .C2 (n_0_0_20));
NOR2_X1 i_0_0_120 (.ZN (n_0_0_50), .A1 (n_0_0_49), .A2 (\i[4] ));
OAI22_X1 i_0_0_119 (.ZN (n_0_0_49), .A1 (n_0_0_14), .A2 (\read_data[10] ), .B1 (\read_data[2] ), .B2 (\i[3] ));
AOI221_X1 i_0_0_118 (.ZN (n_0_0_48), .A (n_0_0_25), .B1 (n_0_0_20), .B2 (\read_data[22] )
    , .C1 (n_0_0_19), .C2 (\read_data[30] ));
OR3_X1 i_0_0_117 (.ZN (n_0_0_47), .A1 (n_0_0_44), .A2 (\i[1] ), .A3 (n_0_0_46));
INV_X1 i_0_0_116 (.ZN (n_0_0_46), .A (n_0_0_45));
OAI221_X1 i_0_0_115 (.ZN (n_0_0_45), .A (n_0_0_20), .B1 (\read_data[16] ), .B2 (\i[2] )
    , .C1 (n_0_0_25), .C2 (\read_data[20] ));
OAI211_X1 i_0_0_114 (.ZN (n_0_0_44), .A (n_0_0_40), .B (n_0_0_41), .C1 (n_0_0_42), .C2 (n_0_0_43));
OAI21_X1 i_0_0_113 (.ZN (n_0_0_43), .A (n_0_0_26), .B1 (\read_data[0] ), .B2 (\i[3] ));
OAI21_X1 i_0_0_112 (.ZN (n_0_0_42), .A (n_0_0_25), .B1 (n_0_0_14), .B2 (\read_data[8] ));
OAI221_X1 i_0_0_111 (.ZN (n_0_0_41), .A (n_0_0_30), .B1 (\read_data[4] ), .B2 (\i[3] )
    , .C1 (n_0_0_14), .C2 (\read_data[12] ));
OAI221_X1 i_0_0_110 (.ZN (n_0_0_40), .A (n_0_0_19), .B1 (\read_data[24] ), .B2 (\i[2] )
    , .C1 (\read_data[28] ), .C2 (n_0_0_25));
OAI21_X1 i_0_0_109 (.ZN (n_0_0_39), .A (n_0_0_29), .B1 (n_0_0_38), .B2 (n_0_0_18));
OAI221_X1 i_0_0_108 (.ZN (n_0_0_38), .A (n_0_0_31), .B1 (n_0_0_35), .B2 (\i[2] ), .C1 (n_0_0_37), .C2 (n_0_0_25));
AOI221_X1 i_0_0_107 (.ZN (n_0_0_37), .A (n_0_0_36), .B1 (\read_data[21] ), .B2 (n_0_0_20)
    , .C1 (\read_data[29] ), .C2 (n_0_0_19));
AND3_X1 i_0_0_106 (.ZN (n_0_0_36), .A1 (n_0_0_26), .A2 (\read_data[13] ), .A3 (\i[3] ));
INV_X1 i_0_0_105 (.ZN (n_0_0_35), .A (n_0_0_34));
OAI21_X1 i_0_0_104 (.ZN (n_0_0_34), .A (n_0_0_32), .B1 (\i[4] ), .B2 (n_0_0_33));
OAI22_X1 i_0_0_103 (.ZN (n_0_0_33), .A1 (n_0_0_14), .A2 (\read_data[9] ), .B1 (\read_data[1] ), .B2 (\i[3] ));
AOI22_X1 i_0_0_102 (.ZN (n_0_0_32), .A1 (\read_data[25] ), .A2 (n_0_0_19), .B1 (n_0_0_20), .B2 (\read_data[17] ));
NAND3_X1 i_0_0_101 (.ZN (n_0_0_31), .A1 (n_0_0_30), .A2 (\read_data[5] ), .A3 (n_0_0_14));
NOR2_X1 i_0_0_100 (.ZN (n_0_0_30), .A1 (n_0_0_25), .A2 (\i[4] ));
OAI221_X1 i_0_0_99 (.ZN (n_0_0_29), .A (n_0_0_18), .B1 (n_0_0_24), .B2 (n_0_0_25)
    , .C1 (n_0_0_28), .C2 (\i[2] ));
AOI221_X1 i_0_0_98 (.ZN (n_0_0_28), .A (n_0_0_27), .B1 (n_0_0_19), .B2 (\read_data[23] )
    , .C1 (\read_data[15] ), .C2 (n_0_0_20));
AND3_X1 i_0_0_97 (.ZN (n_0_0_27), .A1 (n_0_0_26), .A2 (\i[3] ), .A3 (\read_data[7] ));
INV_X1 i_0_0_96 (.ZN (n_0_0_26), .A (\i[4] ));
INV_X1 i_0_0_95 (.ZN (n_0_0_25), .A (\i[2] ));
INV_X1 i_0_0_94 (.ZN (n_0_0_24), .A (n_0_0_23));
OAI21_X1 i_0_0_93 (.ZN (n_0_0_23), .A (n_0_0_21), .B1 (\i[4] ), .B2 (n_0_0_22));
OAI22_X1 i_0_0_92 (.ZN (n_0_0_22), .A1 (n_0_0_14), .A2 (\read_data[11] ), .B1 (\read_data[3] ), .B2 (\i[3] ));
AOI22_X1 i_0_0_91 (.ZN (n_0_0_21), .A1 (n_0_0_19), .A2 (\read_data[27] ), .B1 (n_0_0_20), .B2 (\read_data[19] ));
INV_X1 i_0_0_90 (.ZN (n_0_0_20), .A (n_0_0_15));
INV_X1 i_0_0_89 (.ZN (n_0_0_19), .A (n_0_0_12));
INV_X1 i_0_0_88 (.ZN (n_0_0_18), .A (\i[1] ));
NAND2_X1 i_0_0_87 (.ZN (n_0_131), .A1 (n_0_0_17), .A2 (n_0_0_0));
NOR4_X1 i_0_0_86 (.ZN (n_0_0_17), .A1 (n_0_0_15), .A2 (n_0_0_16), .A3 (\i[2] ), .A4 (\i[1] ));
INV_X1 i_0_0_85 (.ZN (n_0_0_16), .A (\i[0] ));
NAND2_X1 i_0_0_84 (.ZN (n_0_0_15), .A1 (n_0_0_14), .A2 (\i[4] ));
INV_X1 i_0_0_83 (.ZN (n_0_0_14), .A (\i[3] ));
OAI21_X1 i_0_0_82 (.ZN (n_0_130), .A (n_0_0_10), .B1 (n_0_0_13), .B2 (start));
OAI22_X1 i_0_0_81 (.ZN (n_0_0_13), .A1 (n_0_0_11), .A2 (\i[4] ), .B1 (n_0_0_5), .B2 (n_0_0_12));
NAND2_X1 i_0_0_80 (.ZN (n_0_0_12), .A1 (\i[4] ), .A2 (\i[3] ));
INV_X1 i_0_0_79 (.ZN (n_0_0_11), .A (n_0_0_7));
NAND2_X1 i_0_0_78 (.ZN (n_0_0_10), .A1 (start_i[4]), .A2 (start));
NAND2_X1 i_0_0_77 (.ZN (n_0_129), .A1 (n_0_0_8), .A2 (n_0_0_9));
NAND2_X1 i_0_0_76 (.ZN (n_0_0_9), .A1 (start_i[3]), .A2 (start));
OAI211_X1 i_0_0_75 (.ZN (n_0_0_8), .A (n_0_0_7), .B (n_0_0_0), .C1 (\i[3] ), .C2 (n_0_0_6));
NAND2_X1 i_0_0_74 (.ZN (n_0_0_7), .A1 (n_0_0_6), .A2 (\i[3] ));
OAI21_X1 i_0_0_73 (.ZN (n_0_128), .A (n_0_0_3), .B1 (n_0_0_4), .B2 (n_0_0_6));
INV_X1 i_0_0_72 (.ZN (n_0_0_6), .A (n_0_0_5));
NAND2_X1 i_0_0_71 (.ZN (n_0_0_5), .A1 (\i[2] ), .A2 (\i[1] ));
OAI21_X1 i_0_0_70 (.ZN (n_0_0_4), .A (n_0_0_0), .B1 (\i[2] ), .B2 (\i[1] ));
NAND2_X1 i_0_0_69 (.ZN (n_0_0_3), .A1 (start_i[2]), .A2 (start));
AOI22_X1 i_0_0_68 (.ZN (n_0_127), .A1 (n_0_0_2), .A2 (start), .B1 (n_0_0_0), .B2 (\i[1] ));
INV_X1 i_0_0_67 (.ZN (n_0_0_2), .A (start_i[1]));
INV_X1 i_0_0_66 (.ZN (n_0_126), .A (n_0_0_1));
OAI22_X1 i_0_0_65 (.ZN (n_0_0_1), .A1 (n_0_0_0), .A2 (start_i[0]), .B1 (\i[0] ), .B2 (start));
AND2_X1 i_0_0_64 (.ZN (n_0_125), .A1 (n_0_0_0), .A2 (\res[63] ));
AND2_X1 i_0_0_63 (.ZN (n_0_124), .A1 (n_0_0_0), .A2 (\res[62] ));
AND2_X1 i_0_0_62 (.ZN (n_0_123), .A1 (n_0_0_0), .A2 (\res[61] ));
AND2_X1 i_0_0_61 (.ZN (n_0_122), .A1 (hfn_ipo_n24), .A2 (\res[60] ));
AND2_X1 i_0_0_60 (.ZN (n_0_121), .A1 (hfn_ipo_n24), .A2 (\res[59] ));
AND2_X1 i_0_0_59 (.ZN (n_0_120), .A1 (hfn_ipo_n24), .A2 (\res[58] ));
AND2_X1 i_0_0_58 (.ZN (n_0_119), .A1 (hfn_ipo_n24), .A2 (\res[57] ));
AND2_X1 i_0_0_57 (.ZN (n_0_118), .A1 (hfn_ipo_n24), .A2 (\res[56] ));
AND2_X1 i_0_0_56 (.ZN (n_0_117), .A1 (hfn_ipo_n24), .A2 (\res[55] ));
AND2_X1 i_0_0_55 (.ZN (n_0_116), .A1 (hfn_ipo_n24), .A2 (\res[54] ));
AND2_X1 i_0_0_54 (.ZN (n_0_115), .A1 (hfn_ipo_n24), .A2 (\res[53] ));
AND2_X1 i_0_0_53 (.ZN (n_0_114), .A1 (hfn_ipo_n24), .A2 (\res[52] ));
AND2_X1 i_0_0_52 (.ZN (n_0_113), .A1 (hfn_ipo_n24), .A2 (\res[51] ));
AND2_X1 i_0_0_51 (.ZN (n_0_112), .A1 (hfn_ipo_n24), .A2 (\res[50] ));
AND2_X1 i_0_0_50 (.ZN (n_0_111), .A1 (hfn_ipo_n24), .A2 (\res[49] ));
AND2_X1 i_0_0_49 (.ZN (n_0_110), .A1 (hfn_ipo_n24), .A2 (\res[48] ));
AND2_X1 i_0_0_48 (.ZN (n_0_109), .A1 (hfn_ipo_n24), .A2 (\res[47] ));
AND2_X1 i_0_0_47 (.ZN (n_0_108), .A1 (hfn_ipo_n24), .A2 (\res[46] ));
AND2_X1 i_0_0_46 (.ZN (n_0_107), .A1 (hfn_ipo_n24), .A2 (\res[45] ));
AND2_X1 i_0_0_45 (.ZN (n_0_106), .A1 (hfn_ipo_n24), .A2 (\res[44] ));
AND2_X1 i_0_0_44 (.ZN (n_0_105), .A1 (hfn_ipo_n24), .A2 (\res[43] ));
AND2_X1 i_0_0_43 (.ZN (n_0_104), .A1 (hfn_ipo_n24), .A2 (\res[42] ));
AND2_X1 i_0_0_42 (.ZN (n_0_103), .A1 (hfn_ipo_n24), .A2 (\res[41] ));
AND2_X1 i_0_0_41 (.ZN (n_0_102), .A1 (hfn_ipo_n24), .A2 (\res[40] ));
AND2_X1 i_0_0_40 (.ZN (n_0_101), .A1 (hfn_ipo_n24), .A2 (\res[39] ));
AND2_X1 i_0_0_39 (.ZN (n_0_100), .A1 (hfn_ipo_n24), .A2 (\res[38] ));
AND2_X1 i_0_0_38 (.ZN (n_0_99), .A1 (hfn_ipo_n24), .A2 (\res[37] ));
AND2_X1 i_0_0_37 (.ZN (n_0_98), .A1 (hfn_ipo_n24), .A2 (\res[36] ));
AND2_X1 i_0_0_36 (.ZN (n_0_97), .A1 (hfn_ipo_n24), .A2 (\res[35] ));
AND2_X1 i_0_0_35 (.ZN (n_0_96), .A1 (hfn_ipo_n24), .A2 (\res[34] ));
AND2_X1 i_0_0_34 (.ZN (n_0_95), .A1 (hfn_ipo_n24), .A2 (\res[33] ));
AND2_X1 i_0_0_33 (.ZN (n_0_94), .A1 (hfn_ipo_n24), .A2 (\res[32] ));
AND2_X1 i_0_0_32 (.ZN (n_0_93), .A1 (hfn_ipo_n24), .A2 (\res[31] ));
AND2_X1 i_0_0_31 (.ZN (n_0_92), .A1 (hfn_ipo_n24), .A2 (\res[30] ));
AND2_X1 i_0_0_30 (.ZN (n_0_91), .A1 (hfn_ipo_n24), .A2 (\res[29] ));
AND2_X1 i_0_0_29 (.ZN (n_0_90), .A1 (hfn_ipo_n24), .A2 (\res[28] ));
AND2_X1 i_0_0_28 (.ZN (n_0_89), .A1 (hfn_ipo_n24), .A2 (\res[27] ));
AND2_X1 i_0_0_27 (.ZN (n_0_88), .A1 (hfn_ipo_n24), .A2 (\res[26] ));
AND2_X1 i_0_0_26 (.ZN (n_0_87), .A1 (hfn_ipo_n24), .A2 (\res[25] ));
AND2_X1 i_0_0_25 (.ZN (n_0_86), .A1 (hfn_ipo_n24), .A2 (\res[24] ));
AND2_X1 i_0_0_24 (.ZN (n_0_85), .A1 (hfn_ipo_n24), .A2 (\res[23] ));
AND2_X1 i_0_0_23 (.ZN (n_0_84), .A1 (hfn_ipo_n24), .A2 (\res[22] ));
AND2_X1 i_0_0_22 (.ZN (n_0_83), .A1 (hfn_ipo_n24), .A2 (\res[21] ));
AND2_X1 i_0_0_21 (.ZN (n_0_82), .A1 (hfn_ipo_n24), .A2 (\res[20] ));
AND2_X1 i_0_0_20 (.ZN (n_0_81), .A1 (hfn_ipo_n24), .A2 (\res[19] ));
AND2_X1 i_0_0_19 (.ZN (n_0_80), .A1 (hfn_ipo_n24), .A2 (\res[18] ));
AND2_X1 i_0_0_18 (.ZN (n_0_79), .A1 (n_0_0_0), .A2 (\res[17] ));
AND2_X1 i_0_0_17 (.ZN (n_0_78), .A1 (hfn_ipo_n24), .A2 (\res[16] ));
AND2_X1 i_0_0_16 (.ZN (n_0_77), .A1 (hfn_ipo_n24), .A2 (\res[15] ));
AND2_X1 i_0_0_15 (.ZN (n_0_76), .A1 (n_0_0_0), .A2 (\res[14] ));
AND2_X1 i_0_0_14 (.ZN (n_0_75), .A1 (n_0_0_0), .A2 (\res[13] ));
AND2_X1 i_0_0_13 (.ZN (n_0_74), .A1 (n_0_0_0), .A2 (\res[12] ));
AND2_X1 i_0_0_12 (.ZN (n_0_73), .A1 (n_0_0_0), .A2 (\res[11] ));
AND2_X1 i_0_0_11 (.ZN (n_0_72), .A1 (n_0_0_0), .A2 (\res[10] ));
AND2_X1 i_0_0_10 (.ZN (n_0_71), .A1 (n_0_0_0), .A2 (\res[9] ));
AND2_X1 i_0_0_9 (.ZN (n_0_8), .A1 (n_0_0_0), .A2 (\res[8] ));
AND2_X1 i_0_0_8 (.ZN (n_0_7), .A1 (n_0_0_0), .A2 (\res[7] ));
AND2_X1 i_0_0_7 (.ZN (n_0_6), .A1 (n_0_0_0), .A2 (\res[6] ));
AND2_X1 i_0_0_6 (.ZN (n_0_5), .A1 (n_0_0_0), .A2 (\res[5] ));
AND2_X1 i_0_0_5 (.ZN (n_0_4), .A1 (n_0_0_0), .A2 (\res[4] ));
AND2_X1 i_0_0_4 (.ZN (n_0_3), .A1 (n_0_0_0), .A2 (\res[3] ));
AND2_X1 i_0_0_3 (.ZN (n_0_2), .A1 (n_0_0_0), .A2 (\res[2] ));
AND2_X1 i_0_0_2 (.ZN (n_0_1), .A1 (n_0_0_0), .A2 (\res[1] ));
AND2_X1 i_0_0_1 (.ZN (n_0_0), .A1 (n_0_0_0), .A2 (\res[0] ));
INV_X1 i_0_0_0 (.ZN (n_0_0_0), .A (start));
datapath__0_195 i_0_3 (.p_0 ({uc_1, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, 
    n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
    n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
    n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, uc_2}), .p_1 ({1'b0 , \read_data2[31] , 
    \read_data2[30] , \read_data2[29] , \read_data2[28] , \read_data2[27] , \read_data2[26] , 
    \read_data2[25] , \read_data2[24] , \read_data2[23] , \read_data2[22] , \read_data2[21] , 
    \read_data2[20] , \read_data2[19] , \read_data2[18] , \read_data2[17] , \read_data2[16] , 
    \read_data2[15] , \read_data2[14] , \read_data2[13] , \read_data2[12] , \read_data2[11] , 
    \read_data2[10] , \read_data2[9] , \read_data2[8] , \read_data2[7] , \read_data2[6] , 
    \read_data2[5] , \read_data2[4] , \read_data2[3] , \read_data2[2] , \read_data2[1] , 
    \read_data2[0] }));
datapath__0_193 i_0_2 (.p_0 ({n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
    n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, 
    n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
    n_0_12, n_0_11, n_0_10, n_0_9, uc_0}), .read_data2 ({\read_data2[31] , \read_data2[30] , 
    \read_data2[29] , \read_data2[28] , \read_data2[27] , \read_data2[26] , \read_data2[25] , 
    \read_data2[24] , \read_data2[23] , \read_data2[22] , \read_data2[21] , \read_data2[20] , 
    \read_data2[19] , \read_data2[18] , \read_data2[17] , \read_data2[16] , \read_data2[15] , 
    \read_data2[14] , \read_data2[13] , \read_data2[12] , \read_data2[11] , \read_data2[10] , 
    \read_data2[9] , \read_data2[8] , \read_data2[7] , \read_data2[6] , \read_data2[5] , 
    \read_data2[4] , \read_data2[3] , \read_data2[2] , \read_data2[1] , \read_data2[0] }));
DFF_X1 \sum_reg[0]  (.Q (\sum[0] ), .CK (CTS_n_tid1_74), .D (n_0_176));
DFF_X1 \sum_reg[1]  (.Q (\sum[1] ), .CK (CTS_n_tid1_74), .D (n_0_177));
DFF_X1 \sum_reg[2]  (.Q (\sum[2] ), .CK (CTS_n_tid1_74), .D (n_0_178));
DFF_X1 \sum_reg[3]  (.Q (\sum[3] ), .CK (CTS_n_tid1_74), .D (n_0_179));
DFF_X1 \sum_reg[4]  (.Q (\sum[4] ), .CK (CTS_n_tid1_74), .D (n_0_180));
DFF_X1 \sum_reg[5]  (.Q (\sum[5] ), .CK (CTS_n_tid1_74), .D (n_0_181));
DFF_X1 \sum_reg[6]  (.Q (\sum[6] ), .CK (CTS_n_tid1_74), .D (n_0_182));
DFF_X1 \sum_reg[7]  (.Q (\sum[7] ), .CK (CTS_n_tid1_74), .D (n_0_183));
DFF_X1 \sum_reg[8]  (.Q (\sum[8] ), .CK (CTS_n_tid1_74), .D (n_0_184));
DFF_X1 \sum_reg[9]  (.Q (\sum[9] ), .CK (CTS_n_tid1_74), .D (n_0_185));
DFF_X1 \sum_reg[10]  (.Q (\sum[10] ), .CK (CTS_n_tid1_74), .D (n_0_186));
DFF_X1 \sum_reg[11]  (.Q (\sum[11] ), .CK (CTS_n_tid1_74), .D (n_0_187));
DFF_X1 \sum_reg[12]  (.Q (\sum[12] ), .CK (CTS_n_tid1_74), .D (n_0_188));
DFF_X1 \sum_reg[13]  (.Q (\sum[13] ), .CK (CTS_n_tid1_74), .D (n_0_189));
DFF_X1 \sum_reg[14]  (.Q (\sum[14] ), .CK (CTS_n_tid1_74), .D (n_0_190));
DFF_X1 \sum_reg[15]  (.Q (\sum[15] ), .CK (CTS_n_tid1_74), .D (n_0_191));
DFF_X1 \sum_reg[16]  (.Q (\sum[16] ), .CK (CTS_n_tid1_74), .D (n_0_192));
DFF_X1 \sum_reg[17]  (.Q (\sum[17] ), .CK (CTS_n_tid1_74), .D (n_0_193));
DFF_X1 \sum_reg[18]  (.Q (\sum[18] ), .CK (CTS_n_tid1_75), .D (n_0_194));
DFF_X1 \sum_reg[19]  (.Q (\sum[19] ), .CK (CTS_n_tid1_75), .D (n_0_195));
DFF_X1 \sum_reg[20]  (.Q (\sum[20] ), .CK (CTS_n_tid1_75), .D (n_0_196));
DFF_X1 \sum_reg[21]  (.Q (\sum[21] ), .CK (CTS_n_tid1_75), .D (n_0_197));
DFF_X1 \sum_reg[22]  (.Q (\sum[22] ), .CK (CTS_n_tid1_75), .D (n_0_198));
DFF_X1 \sum_reg[23]  (.Q (\sum[23] ), .CK (CTS_n_tid1_75), .D (n_0_199));
DFF_X1 \sum_reg[24]  (.Q (\sum[24] ), .CK (CTS_n_tid1_75), .D (n_0_200));
DFF_X1 \sum_reg[25]  (.Q (\sum[25] ), .CK (CTS_n_tid1_75), .D (n_0_201));
DFF_X1 \sum_reg[26]  (.Q (\sum[26] ), .CK (CTS_n_tid1_75), .D (n_0_132));
DFF_X1 \sum_reg[27]  (.Q (\sum[27] ), .CK (CTS_n_tid1_75), .D (n_0_133));
DFF_X1 \sum_reg[28]  (.Q (\sum[28] ), .CK (CTS_n_tid1_75), .D (n_0_134));
DFF_X1 \sum_reg[29]  (.Q (\sum[29] ), .CK (CTS_n_tid1_75), .D (n_0_135));
DFF_X1 \sum_reg[30]  (.Q (\sum[30] ), .CK (CTS_n_tid1_75), .D (n_0_136));
DFF_X1 \sum_reg[31]  (.Q (\sum[31] ), .CK (CTS_n_tid1_75), .D (n_0_137));
DFF_X1 \sum_reg[32]  (.Q (\sum[32] ), .CK (CTS_n_tid1_75), .D (n_0_138));
DFF_X1 \sum_reg[33]  (.Q (\sum[33] ), .CK (CTS_n_tid1_75), .D (n_0_139));
DFF_X1 \sum_reg[34]  (.Q (\sum[34] ), .CK (CTS_n_tid1_75), .D (n_0_140));
DFF_X1 \sum_reg[35]  (.Q (\sum[35] ), .CK (CTS_n_tid1_75), .D (n_0_141));
DFF_X1 \sum_reg[36]  (.Q (\sum[36] ), .CK (CTS_n_tid1_75), .D (n_0_142));
DFF_X1 \sum_reg[37]  (.Q (\sum[37] ), .CK (CTS_n_tid1_75), .D (n_0_143));
DFF_X1 \sum_reg[38]  (.Q (\sum[38] ), .CK (CTS_n_tid1_55), .D (n_0_144));
DFF_X1 \sum_reg[39]  (.Q (\sum[39] ), .CK (CTS_n_tid1_75), .D (n_0_145));
DFF_X1 \sum_reg[40]  (.Q (\sum[40] ), .CK (CTS_n_tid1_55), .D (n_0_146));
DFF_X1 \sum_reg[41]  (.Q (\sum[41] ), .CK (CTS_n_tid1_55), .D (n_0_147));
DFF_X1 \sum_reg[42]  (.Q (\sum[42] ), .CK (CTS_n_tid1_55), .D (n_0_148));
DFF_X1 \sum_reg[43]  (.Q (\sum[43] ), .CK (CTS_n_tid1_55), .D (n_0_149));
DFF_X1 \sum_reg[44]  (.Q (\sum[44] ), .CK (CTS_n_tid1_55), .D (n_0_150));
DFF_X1 \sum_reg[45]  (.Q (\sum[45] ), .CK (CTS_n_tid1_55), .D (n_0_151));
DFF_X1 \sum_reg[46]  (.Q (\sum[46] ), .CK (CTS_n_tid1_55), .D (n_0_152));
DFF_X1 \sum_reg[47]  (.Q (\sum[47] ), .CK (CTS_n_tid1_55), .D (n_0_153));
DFF_X1 \sum_reg[48]  (.Q (\sum[48] ), .CK (CTS_n_tid1_55), .D (n_0_154));
DFF_X1 \sum_reg[49]  (.Q (\sum[49] ), .CK (CTS_n_tid1_55), .D (n_0_155));
DFF_X1 \sum_reg[50]  (.Q (\sum[50] ), .CK (CTS_n_tid1_55), .D (n_0_156));
DFF_X1 \sum_reg[51]  (.Q (\sum[51] ), .CK (CTS_n_tid1_55), .D (n_0_157));
DFF_X1 \sum_reg[52]  (.Q (\sum[52] ), .CK (CTS_n_tid1_55), .D (n_0_158));
DFF_X1 \sum_reg[53]  (.Q (\sum[53] ), .CK (CTS_n_tid1_55), .D (n_0_159));
DFF_X1 \sum_reg[54]  (.Q (\sum[54] ), .CK (CTS_n_tid1_55), .D (n_0_160));
DFF_X1 \sum_reg[55]  (.Q (\sum[55] ), .CK (CTS_n_tid1_55), .D (n_0_161));
DFF_X1 \sum_reg[56]  (.Q (\sum[56] ), .CK (CTS_n_tid1_55), .D (n_0_162));
DFF_X1 \sum_reg[57]  (.Q (\sum[57] ), .CK (CTS_n_tid1_55), .D (n_0_163));
DFF_X1 \sum_reg[58]  (.Q (\sum[58] ), .CK (CTS_n_tid1_55), .D (n_0_164));
DFF_X1 \sum_reg[59]  (.Q (\sum[59] ), .CK (CTS_n_tid1_55), .D (n_0_165));
DFF_X1 \sum_reg[60]  (.Q (\sum[60] ), .CK (CTS_n_tid1_55), .D (n_0_166));
DFF_X1 \sum_reg[61]  (.Q (\sum[61] ), .CK (CTS_n_tid1_55), .D (n_0_167));
DFF_X1 \sum_reg[62]  (.Q (\sum[62] ), .CK (CTS_n_tid1_55), .D (n_0_168));
DFF_X1 \sum_reg[63]  (.Q (\sum[63] ), .CK (CTS_n_tid1_55), .D (n_0_169));
regFile64 r2 (.read_data ({read_data3[63], read_data3[62], read_data3[61], read_data3[60], 
    read_data3[59], read_data3[58], read_data3[57], read_data3[56], read_data3[55], 
    read_data3[54], read_data3[53], read_data3[52], read_data3[51], read_data3[50], 
    read_data3[49], read_data3[48], read_data3[47], read_data3[46], read_data3[45], 
    read_data3[44], read_data3[43], read_data3[42], read_data3[41], read_data3[40], 
    read_data3[39], read_data3[38], read_data3[37], read_data3[36], read_data3[35], 
    read_data3[34], read_data3[33], read_data3[32], read_data3[31], read_data3[30], 
    read_data3[29], read_data3[28], read_data3[27], read_data3[26], read_data3[25], 
    read_data3[24], read_data3[23], read_data3[22], read_data3[21], read_data3[20], 
    read_data3[19], read_data3[18], read_data3[17], read_data3[16], read_data3[15], 
    read_data3[14], read_data3[13], read_data3[12], read_data3[11], read_data3[10], 
    read_data3[9], read_data3[8], read_data3[7], read_data3[6], read_data3[5], read_data3[4], 
    read_data3[3], read_data3[2], read_data3[1], read_data3[0]}), .write_data ({\res[63] , 
    \res[62] , \res[61] , \res[60] , \res[59] , \res[58] , \res[57] , \res[56] , 
    \res[55] , \res[54] , \res[53] , \res[52] , \res[51] , \res[50] , \res[49] , 
    \res[48] , \res[47] , \res[46] , \res[45] , \res[44] , \res[43] , \res[42] , 
    \res[41] , \res[40] , \res[39] , \res[38] , \res[37] , \res[36] , \res[35] , 
    \res[34] , \res[33] , \res[32] , \res[31] , \res[30] , \res[29] , \res[28] , 
    \res[27] , \res[26] , \res[25] , \res[24] , \res[23] , \res[22] , \res[21] , 
    \res[20] , \res[19] , \res[18] , \res[17] , \res[16] , \res[15] , \res[14] , 
    \res[13] , \res[12] , \res[11] , \res[10] , \res[9] , \res[8] , \res[7] , \res[6] , 
    \res[5] , \res[4] , \res[3] , \res[2] , \res[1] , \res[0] }), .clk__CTS_1_PP_1 (n_tid1_110));
carry_lookahead_adder ADD (.o_result ({\res[63] , \res[62] , \res[61] , \res[60] , 
    \res[59] , \res[58] , \res[57] , \res[56] , \res[55] , \res[54] , \res[53] , 
    \res[52] , \res[51] , \res[50] , \res[49] , \res[48] , \res[47] , \res[46] , 
    \res[45] , \res[44] , \res[43] , \res[42] , \res[41] , \res[40] , \res[39] , 
    \res[38] , \res[37] , \res[36] , \res[35] , \res[34] , \res[33] , \res[32] , 
    \res[31] , \res[30] , \res[29] , \res[28] , \res[27] , \res[26] , \res[25] , 
    \res[24] , \res[23] , \res[22] , \res[21] , \res[20] , \res[19] , \res[18] , 
    \res[17] , \res[16] , \res[15] , \res[14] , \res[13] , \res[12] , \res[11] , 
    \res[10] , \res[9] , \res[8] , \res[7] , \res[6] , \res[5] , \res[4] , \res[3] , 
    \res[2] , \res[1] , \res[0] }), .i_add1 ({\c[63] , \c[62] , \c[61] , \c[60] , 
    \c[59] , \c[58] , \c[57] , \c[56] , \c[55] , \c[54] , \c[53] , \c[52] , \c[51] , 
    \c[50] , \c[49] , \c[48] , \c[47] , \c[46] , \c[45] , \c[44] , \c[43] , \c[42] , 
    \c[41] , \c[40] , \c[39] , \c[38] , \c[37] , \c[36] , \c[35] , \c[34] , \c[33] , 
    \c[32] , \c[31] , \c[30] , \c[29] , \c[28] , \c[27] , \c[26] , \c[25] , \c[24] , 
    \c[23] , \c[22] , \c[21] , \c[20] , \c[19] , \c[18] , \c[17] , \c[16] , \c[15] , 
    \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , \c[8] , \c[7] , \c[6] , 
    \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] }), .i_add2 ({\sum[63] , \sum[62] , 
    \sum[61] , \sum[60] , \sum[59] , \sum[58] , \sum[57] , \sum[56] , \sum[55] , 
    \sum[54] , \sum[53] , \sum[52] , \sum[51] , \sum[50] , \sum[49] , \sum[48] , 
    \sum[47] , \sum[46] , \sum[45] , \sum[44] , \sum[43] , \sum[42] , \sum[41] , 
    \sum[40] , \sum[39] , \sum[38] , \sum[37] , \sum[36] , \sum[35] , \sum[34] , 
    \sum[33] , \sum[32] , \sum[31] , \sum[30] , \sum[29] , \sum[28] , \sum[27] , 
    \sum[26] , \sum[25] , \sum[24] , \sum[23] , \sum[22] , \sum[21] , \sum[20] , 
    \sum[19] , \sum[18] , \sum[17] , \sum[16] , \sum[15] , \sum[14] , \sum[13] , 
    \sum[12] , \sum[11] , \sum[10] , \sum[9] , \sum[8] , \sum[7] , \sum[6] , \sum[5] , 
    \sum[4] , \sum[3] , \sum[2] , \sum[1] , \sum[0] }));
regFile r (.read_data2 ({\read_data2[31] , \read_data2[30] , \read_data2[29] , \read_data2[28] , 
    \read_data2[27] , \read_data2[26] , \read_data2[25] , \read_data2[24] , \read_data2[23] , 
    \read_data2[22] , \read_data2[21] , \read_data2[20] , \read_data2[19] , \read_data2[18] , 
    \read_data2[17] , \read_data2[16] , \read_data2[15] , \read_data2[14] , \read_data2[13] , 
    \read_data2[12] , \read_data2[11] , \read_data2[10] , \read_data2[9] , \read_data2[8] , 
    \read_data2[7] , \read_data2[6] , \read_data2[5] , \read_data2[4] , \read_data2[3] , 
    \read_data2[2] , \read_data2[1] , \read_data2[0] }), .read_data ({\read_data[31] , 
    \read_data[30] , \read_data[29] , \read_data[28] , \read_data[27] , \read_data[26] , 
    \read_data[25] , \read_data[24] , \read_data[23] , \read_data[22] , \read_data[21] , 
    \read_data[20] , \read_data[19] , \read_data[18] , \read_data[17] , \read_data[16] , 
    \read_data[15] , \read_data[14] , \read_data[13] , \read_data[12] , \read_data[11] , 
    \read_data[10] , \read_data[9] , \read_data[8] , \read_data[7] , \read_data[6] , 
    \read_data[5] , \read_data[4] , \read_data[3] , \read_data[2] , \read_data[1] , 
    \read_data[0] }), .write_data2 ({b[31], b[30], b[29], b[28], b[27], b[26], b[25], 
    b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], b[15], b[14], 
    b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], 
    b[0]}), .write_data ({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24], 
    a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], a[13], 
    a[12], a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]})
    , .write_en (write_en), .clk__CTS_1_PP_1 (n_tid1_110));
CLKBUF_X3 CTS_L1_tid1__c1_tid1__c85 (.Z (n_tid1_110), .A (clk));
BUF_X2 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (n_0_0_0));
CLKBUF_X1 hfn_ipo_c32 (.Z (hfn_ipo_n32), .A (\shift[1] ));
BUF_X4 drc_ipo_c33 (.Z (drc_ipo_n33), .A (\shift[2] ));
CLKBUF_X1 hfn_ipo_c25 (.Z (hfn_ipo_n25), .A (n_0_0_101));
CLKBUF_X2 CTS_L2_c_tid1_77 (.Z (CTS_n_tid1_74), .A (n_tid1_110));
CLKBUF_X1 hfn_ipo_c27 (.Z (hfn_ipo_n27), .A (n_0_0_108));
CLKBUF_X2 CTS_L2_c_tid1_58 (.Z (CTS_n_tid1_55), .A (n_tid1_110));
CLKBUF_X1 hfn_ipo_c31 (.Z (hfn_ipo_n31), .A (\shift[1] ));
CLKBUF_X1 hfn_ipo_c29 (.Z (hfn_ipo_n29), .A (n_0_0_109));
BUF_X4 drc_ipo_c34 (.Z (drc_ipo_n34), .A (\shift[3] ));
CLKBUF_X2 CTS_L2_c_tid1_78 (.Z (CTS_n_tid1_75), .A (n_tid1_110));

endmodule //Radix4


