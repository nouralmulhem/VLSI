/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 14:15:26 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2616278483 */

module regFile(read_data, read_data2, write_en, write_data, write_data2, clk);
   output [31:0]read_data;
   output [31:0]read_data2;
   input write_en;
   input [31:0]write_data;
   input [31:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[31]  (.D(write_data2[31]), .CK(n_0), .Q(read_data2[31]), 
      .QN());
   DFF_X1 \my_reg2_reg[30]  (.D(write_data2[30]), .CK(n_0), .Q(read_data2[30]), 
      .QN());
   DFF_X1 \my_reg2_reg[29]  (.D(write_data2[29]), .CK(n_0), .Q(read_data2[29]), 
      .QN());
   DFF_X1 \my_reg2_reg[28]  (.D(write_data2[28]), .CK(n_0), .Q(read_data2[28]), 
      .QN());
   DFF_X1 \my_reg2_reg[27]  (.D(write_data2[27]), .CK(n_0), .Q(read_data2[27]), 
      .QN());
   DFF_X1 \my_reg2_reg[26]  (.D(write_data2[26]), .CK(n_0), .Q(read_data2[26]), 
      .QN());
   DFF_X1 \my_reg2_reg[25]  (.D(write_data2[25]), .CK(n_0), .Q(read_data2[25]), 
      .QN());
   DFF_X1 \my_reg2_reg[24]  (.D(write_data2[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data2[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
   DFF_X1 \my_reg2_reg[22]  (.D(write_data2[22]), .CK(n_0), .Q(read_data2[22]), 
      .QN());
   DFF_X1 \my_reg2_reg[21]  (.D(write_data2[21]), .CK(n_0), .Q(read_data2[21]), 
      .QN());
   DFF_X1 \my_reg2_reg[20]  (.D(write_data2[20]), .CK(n_0), .Q(read_data2[20]), 
      .QN());
   DFF_X1 \my_reg2_reg[19]  (.D(write_data2[19]), .CK(n_0), .Q(read_data2[19]), 
      .QN());
   DFF_X1 \my_reg2_reg[18]  (.D(write_data2[18]), .CK(n_0), .Q(read_data2[18]), 
      .QN());
   DFF_X1 \my_reg2_reg[17]  (.D(write_data2[17]), .CK(n_0), .Q(read_data2[17]), 
      .QN());
   DFF_X1 \my_reg2_reg[16]  (.D(write_data2[16]), .CK(n_0), .Q(read_data2[16]), 
      .QN());
   DFF_X1 \my_reg2_reg[15]  (.D(write_data2[15]), .CK(n_0), .Q(read_data2[15]), 
      .QN());
   DFF_X1 \my_reg2_reg[14]  (.D(write_data2[14]), .CK(n_0), .Q(read_data2[14]), 
      .QN());
   DFF_X1 \my_reg2_reg[13]  (.D(write_data2[13]), .CK(n_0), .Q(read_data2[13]), 
      .QN());
   DFF_X1 \my_reg2_reg[12]  (.D(write_data2[12]), .CK(n_0), .Q(read_data2[12]), 
      .QN());
   DFF_X1 \my_reg2_reg[11]  (.D(write_data2[11]), .CK(n_0), .Q(read_data2[11]), 
      .QN());
   DFF_X1 \my_reg2_reg[10]  (.D(write_data2[10]), .CK(n_0), .Q(read_data2[10]), 
      .QN());
   DFF_X1 \my_reg2_reg[9]  (.D(write_data2[9]), .CK(n_0), .Q(read_data2[9]), 
      .QN());
   DFF_X1 \my_reg2_reg[8]  (.D(write_data2[8]), .CK(n_0), .Q(read_data2[8]), 
      .QN());
   DFF_X1 \my_reg2_reg[7]  (.D(write_data2[7]), .CK(n_0), .Q(read_data2[7]), 
      .QN());
   DFF_X1 \my_reg2_reg[6]  (.D(write_data2[6]), .CK(n_0), .Q(read_data2[6]), 
      .QN());
   DFF_X1 \my_reg2_reg[5]  (.D(write_data2[5]), .CK(n_0), .Q(read_data2[5]), 
      .QN());
   DFF_X1 \my_reg2_reg[4]  (.D(write_data2[4]), .CK(n_0), .Q(read_data2[4]), 
      .QN());
   DFF_X1 \my_reg2_reg[3]  (.D(write_data2[3]), .CK(n_0), .Q(read_data2[3]), 
      .QN());
   DFF_X1 \my_reg2_reg[2]  (.D(write_data2[2]), .CK(n_0), .Q(read_data2[2]), 
      .QN());
   DFF_X1 \my_reg2_reg[1]  (.D(write_data2[1]), .CK(n_0), .Q(read_data2[1]), 
      .QN());
   DFF_X1 \my_reg2_reg[0]  (.D(write_data2[0]), .CK(n_0), .Q(read_data2[0]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
endmodule

module regFile64(read_data, write_en, write_data, clk);
   output [63:0]read_data;
   input write_en;
   input [63:0]write_data;
   input clk;

   DFF_X1 \my_reg_reg[63]  (.D(write_data[63]), .CK(n_0), .Q(read_data[63]), 
      .QN());
   INV_X1 i_0_0 (.A(clk), .ZN(n_0));
   DFF_X1 \my_reg_reg[62]  (.D(write_data[62]), .CK(n_0), .Q(read_data[62]), 
      .QN());
   DFF_X1 \my_reg_reg[61]  (.D(write_data[61]), .CK(n_0), .Q(read_data[61]), 
      .QN());
   DFF_X1 \my_reg_reg[60]  (.D(write_data[60]), .CK(n_0), .Q(read_data[60]), 
      .QN());
   DFF_X1 \my_reg_reg[59]  (.D(write_data[59]), .CK(n_0), .Q(read_data[59]), 
      .QN());
   DFF_X1 \my_reg_reg[58]  (.D(write_data[58]), .CK(n_0), .Q(read_data[58]), 
      .QN());
   DFF_X1 \my_reg_reg[57]  (.D(write_data[57]), .CK(n_0), .Q(read_data[57]), 
      .QN());
   DFF_X1 \my_reg_reg[56]  (.D(write_data[56]), .CK(n_0), .Q(read_data[56]), 
      .QN());
   DFF_X1 \my_reg_reg[55]  (.D(write_data[55]), .CK(n_0), .Q(read_data[55]), 
      .QN());
   DFF_X1 \my_reg_reg[54]  (.D(write_data[54]), .CK(n_0), .Q(read_data[54]), 
      .QN());
   DFF_X1 \my_reg_reg[53]  (.D(write_data[53]), .CK(n_0), .Q(read_data[53]), 
      .QN());
   DFF_X1 \my_reg_reg[52]  (.D(write_data[52]), .CK(n_0), .Q(read_data[52]), 
      .QN());
   DFF_X1 \my_reg_reg[51]  (.D(write_data[51]), .CK(n_0), .Q(read_data[51]), 
      .QN());
   DFF_X1 \my_reg_reg[50]  (.D(write_data[50]), .CK(n_0), .Q(read_data[50]), 
      .QN());
   DFF_X1 \my_reg_reg[49]  (.D(write_data[49]), .CK(n_0), .Q(read_data[49]), 
      .QN());
   DFF_X1 \my_reg_reg[48]  (.D(write_data[48]), .CK(n_0), .Q(read_data[48]), 
      .QN());
   DFF_X1 \my_reg_reg[47]  (.D(write_data[47]), .CK(n_0), .Q(read_data[47]), 
      .QN());
   DFF_X1 \my_reg_reg[46]  (.D(write_data[46]), .CK(n_0), .Q(read_data[46]), 
      .QN());
   DFF_X1 \my_reg_reg[45]  (.D(write_data[45]), .CK(n_0), .Q(read_data[45]), 
      .QN());
   DFF_X1 \my_reg_reg[44]  (.D(write_data[44]), .CK(n_0), .Q(read_data[44]), 
      .QN());
   DFF_X1 \my_reg_reg[43]  (.D(write_data[43]), .CK(n_0), .Q(read_data[43]), 
      .QN());
   DFF_X1 \my_reg_reg[42]  (.D(write_data[42]), .CK(n_0), .Q(read_data[42]), 
      .QN());
   DFF_X1 \my_reg_reg[41]  (.D(write_data[41]), .CK(n_0), .Q(read_data[41]), 
      .QN());
   DFF_X1 \my_reg_reg[40]  (.D(write_data[40]), .CK(n_0), .Q(read_data[40]), 
      .QN());
   DFF_X1 \my_reg_reg[39]  (.D(write_data[39]), .CK(n_0), .Q(read_data[39]), 
      .QN());
   DFF_X1 \my_reg_reg[38]  (.D(write_data[38]), .CK(n_0), .Q(read_data[38]), 
      .QN());
   DFF_X1 \my_reg_reg[37]  (.D(write_data[37]), .CK(n_0), .Q(read_data[37]), 
      .QN());
   DFF_X1 \my_reg_reg[36]  (.D(write_data[36]), .CK(n_0), .Q(read_data[36]), 
      .QN());
   DFF_X1 \my_reg_reg[35]  (.D(write_data[35]), .CK(n_0), .Q(read_data[35]), 
      .QN());
   DFF_X1 \my_reg_reg[34]  (.D(write_data[34]), .CK(n_0), .Q(read_data[34]), 
      .QN());
   DFF_X1 \my_reg_reg[33]  (.D(write_data[33]), .CK(n_0), .Q(read_data[33]), 
      .QN());
   DFF_X1 \my_reg_reg[32]  (.D(write_data[32]), .CK(n_0), .Q(read_data[32]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
endmodule

module datapath(p_0, read_data2);
   output [31:0]p_0;
   input [31:0]read_data2;

   XOR2_X1 i_0 (.A(read_data2[1]), .B(read_data2[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(read_data2[2]), .B1(read_data2[1]), .B2(read_data2[0]), 
      .ZN(n_0));
   XOR2_X1 i_3 (.A(read_data2[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(read_data2[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(read_data2[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(read_data2[6]), .B1(n_27), .B2(read_data2[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(read_data2[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(read_data2[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(read_data2[9]), .B1(n_25), .B2(read_data2[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(read_data2[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(read_data2[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(read_data2[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(read_data2[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(read_data2[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(read_data2[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(read_data2[16]), .B1(n_19), .B2(read_data2[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(read_data2[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(read_data2[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(read_data2[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(read_data2[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(read_data2[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(read_data2[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(read_data2[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(read_data2[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(read_data2[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(read_data2[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(read_data2[27]), .B1(n_9), .B2(read_data2[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(read_data2[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(read_data2[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(read_data2[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(read_data2[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(read_data2[28]), .A3(read_data2[29]), .A4(
      read_data2[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(read_data2[28]), .A3(read_data2[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(read_data2[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(read_data2[26]), .A3(read_data2[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(read_data2[23]), .A3(read_data2[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(read_data2[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(read_data2[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(read_data2[18]), .A3(read_data2[19]), .A4(
      read_data2[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(read_data2[18]), .A3(read_data2[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(read_data2[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(read_data2[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(read_data2[15]), .A3(read_data2[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(read_data2[12]), .A3(read_data2[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(read_data2[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(read_data2[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(read_data2[8]), .A3(read_data2[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(read_data2[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(read_data2[5]), .A3(read_data2[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(read_data2[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(read_data2[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(read_data2[2]), .A2(read_data2[1]), .A3(read_data2[0]), 
      .ZN(n_29));
   INV_X1 i_61 (.A(read_data2[11]), .ZN(n_30));
   INV_X1 i_62 (.A(read_data2[14]), .ZN(n_31));
   INV_X1 i_63 (.A(read_data2[21]), .ZN(n_32));
   INV_X1 i_64 (.A(read_data2[25]), .ZN(n_33));
endmodule

module datapath__0_128(p_0, p_1);
   output [32:0]p_0;
   input [32:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_27), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_25), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(p_1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(p_1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(p_1[16]), .B1(n_19), .B2(p_1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(p_1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(p_1[27]), .B1(n_9), .B2(p_1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(p_1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(p_1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(p_1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(p_1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(p_1[26]), .A3(p_1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(p_1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(p_1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(p_1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(p_1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(p_1[15]), .A3(p_1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(p_1[12]), .A3(p_1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(p_1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(p_1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(p_1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(p_1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(p_1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(p_1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(p_1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(p_1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(p_1[25]), .ZN(n_33));
endmodule

module datapath__0_142(c, p_0, p_1);
   input [63:0]c;
   input [63:0]p_0;
   output [63:0]p_1;

   AOI21_X1 i_0 (.A(n_132), .B1(n_200), .B2(n_197), .ZN(p_1[0]));
   XNOR2_X1 i_1 (.A(n_132), .B(n_0), .ZN(p_1[1]));
   OAI22_X1 i_2 (.A1(n_201), .A2(n_198), .B1(c[1]), .B2(p_0[1]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(n_134), .B(n_130), .ZN(p_1[2]));
   XNOR2_X1 i_4 (.A(n_129), .B(n_127), .ZN(p_1[3]));
   XNOR2_X1 i_5 (.A(n_126), .B(n_124), .ZN(p_1[4]));
   XNOR2_X1 i_6 (.A(n_123), .B(n_121), .ZN(p_1[5]));
   XNOR2_X1 i_7 (.A(n_120), .B(n_118), .ZN(p_1[6]));
   XNOR2_X1 i_8 (.A(n_117), .B(n_115), .ZN(p_1[7]));
   XNOR2_X1 i_9 (.A(n_114), .B(n_112), .ZN(p_1[8]));
   XNOR2_X1 i_10 (.A(n_111), .B(n_109), .ZN(p_1[9]));
   XNOR2_X1 i_11 (.A(n_108), .B(n_106), .ZN(p_1[10]));
   XNOR2_X1 i_12 (.A(n_105), .B(n_103), .ZN(p_1[11]));
   XNOR2_X1 i_13 (.A(n_102), .B(n_100), .ZN(p_1[12]));
   XNOR2_X1 i_14 (.A(n_99), .B(n_97), .ZN(p_1[13]));
   XNOR2_X1 i_15 (.A(n_96), .B(n_94), .ZN(p_1[14]));
   XOR2_X1 i_16 (.A(n_93), .B(n_92), .Z(p_1[15]));
   XNOR2_X1 i_17 (.A(n_91), .B(n_1), .ZN(p_1[16]));
   OAI22_X1 i_18 (.A1(c[16]), .A2(p_0[16]), .B1(n_202), .B2(n_199), .ZN(n_1));
   XNOR2_X1 i_19 (.A(n_137), .B(n_89), .ZN(p_1[17]));
   XNOR2_X1 i_20 (.A(n_88), .B(n_86), .ZN(p_1[18]));
   XNOR2_X1 i_21 (.A(n_85), .B(n_83), .ZN(p_1[19]));
   XNOR2_X1 i_22 (.A(n_82), .B(n_80), .ZN(p_1[20]));
   XOR2_X1 i_23 (.A(n_79), .B(n_2), .Z(p_1[21]));
   OAI21_X1 i_24 (.A(n_139), .B1(c[21]), .B2(p_0[21]), .ZN(n_2));
   XNOR2_X1 i_25 (.A(n_141), .B(n_78), .ZN(p_1[22]));
   XOR2_X1 i_26 (.A(n_77), .B(n_3), .Z(p_1[23]));
   OAI21_X1 i_27 (.A(n_142), .B1(c[23]), .B2(p_0[23]), .ZN(n_3));
   XOR2_X1 i_28 (.A(n_143), .B(n_75), .Z(p_1[24]));
   XOR2_X1 i_29 (.A(n_74), .B(n_73), .Z(p_1[25]));
   XOR2_X1 i_30 (.A(n_72), .B(n_4), .Z(p_1[26]));
   OAI21_X1 i_31 (.A(n_146), .B1(c[26]), .B2(p_0[26]), .ZN(n_4));
   XNOR2_X1 i_32 (.A(n_148), .B(n_71), .ZN(p_1[27]));
   XOR2_X1 i_33 (.A(n_70), .B(n_5), .Z(p_1[28]));
   OAI21_X1 i_34 (.A(n_149), .B1(c[28]), .B2(p_0[28]), .ZN(n_5));
   XOR2_X1 i_35 (.A(n_150), .B(n_68), .Z(p_1[29]));
   XOR2_X1 i_36 (.A(n_67), .B(n_66), .Z(p_1[30]));
   XOR2_X1 i_37 (.A(n_65), .B(n_6), .Z(p_1[31]));
   OAI21_X1 i_38 (.A(n_153), .B1(c[31]), .B2(p_0[31]), .ZN(n_6));
   XNOR2_X1 i_39 (.A(n_155), .B(n_64), .ZN(p_1[32]));
   XOR2_X1 i_40 (.A(n_63), .B(n_7), .Z(p_1[33]));
   OAI21_X1 i_41 (.A(n_156), .B1(c[33]), .B2(p_0[33]), .ZN(n_7));
   XOR2_X1 i_42 (.A(n_157), .B(n_61), .Z(p_1[34]));
   XOR2_X1 i_43 (.A(n_60), .B(n_59), .Z(p_1[35]));
   XOR2_X1 i_44 (.A(n_58), .B(n_8), .Z(p_1[36]));
   OAI21_X1 i_45 (.A(n_160), .B1(c[36]), .B2(p_0[36]), .ZN(n_8));
   XNOR2_X1 i_46 (.A(n_162), .B(n_57), .ZN(p_1[37]));
   XOR2_X1 i_47 (.A(n_56), .B(n_9), .Z(p_1[38]));
   OAI21_X1 i_48 (.A(n_163), .B1(c[38]), .B2(p_0[38]), .ZN(n_9));
   XOR2_X1 i_49 (.A(n_164), .B(n_54), .Z(p_1[39]));
   XOR2_X1 i_50 (.A(n_53), .B(n_52), .Z(p_1[40]));
   XOR2_X1 i_51 (.A(n_51), .B(n_10), .Z(p_1[41]));
   OAI21_X1 i_52 (.A(n_167), .B1(c[41]), .B2(p_0[41]), .ZN(n_10));
   XNOR2_X1 i_53 (.A(n_169), .B(n_50), .ZN(p_1[42]));
   XOR2_X1 i_54 (.A(n_49), .B(n_11), .Z(p_1[43]));
   OAI21_X1 i_55 (.A(n_170), .B1(c[43]), .B2(p_0[43]), .ZN(n_11));
   XOR2_X1 i_56 (.A(n_171), .B(n_47), .Z(p_1[44]));
   XOR2_X1 i_57 (.A(n_46), .B(n_45), .Z(p_1[45]));
   XOR2_X1 i_58 (.A(n_44), .B(n_12), .Z(p_1[46]));
   OAI21_X1 i_59 (.A(n_174), .B1(c[46]), .B2(p_0[46]), .ZN(n_12));
   XNOR2_X1 i_60 (.A(n_176), .B(n_43), .ZN(p_1[47]));
   XOR2_X1 i_61 (.A(n_42), .B(n_13), .Z(p_1[48]));
   OAI21_X1 i_62 (.A(n_177), .B1(c[48]), .B2(p_0[48]), .ZN(n_13));
   XOR2_X1 i_63 (.A(n_178), .B(n_40), .Z(p_1[49]));
   XOR2_X1 i_64 (.A(n_39), .B(n_38), .Z(p_1[50]));
   XOR2_X1 i_65 (.A(n_37), .B(n_14), .Z(p_1[51]));
   OAI21_X1 i_66 (.A(n_181), .B1(c[51]), .B2(p_0[51]), .ZN(n_14));
   XNOR2_X1 i_67 (.A(n_183), .B(n_36), .ZN(p_1[52]));
   XOR2_X1 i_68 (.A(n_35), .B(n_15), .Z(p_1[53]));
   OAI21_X1 i_69 (.A(n_184), .B1(c[53]), .B2(p_0[53]), .ZN(n_15));
   XOR2_X1 i_70 (.A(n_185), .B(n_33), .Z(p_1[54]));
   XOR2_X1 i_71 (.A(n_32), .B(n_31), .Z(p_1[55]));
   XOR2_X1 i_72 (.A(n_30), .B(n_16), .Z(p_1[56]));
   OAI21_X1 i_73 (.A(n_188), .B1(c[56]), .B2(p_0[56]), .ZN(n_16));
   XNOR2_X1 i_74 (.A(n_190), .B(n_29), .ZN(p_1[57]));
   XOR2_X1 i_75 (.A(n_28), .B(n_17), .Z(p_1[58]));
   OAI21_X1 i_76 (.A(n_191), .B1(c[58]), .B2(p_0[58]), .ZN(n_17));
   XOR2_X1 i_77 (.A(n_192), .B(n_26), .Z(p_1[59]));
   XOR2_X1 i_78 (.A(n_25), .B(n_24), .Z(p_1[60]));
   XOR2_X1 i_79 (.A(n_23), .B(n_18), .Z(p_1[61]));
   OAI21_X1 i_80 (.A(n_194), .B1(c[61]), .B2(p_0[61]), .ZN(n_18));
   XOR2_X1 i_81 (.A(n_195), .B(n_21), .Z(p_1[62]));
   XOR2_X1 i_82 (.A(n_20), .B(n_19), .Z(p_1[63]));
   XOR2_X1 i_83 (.A(c[63]), .B(p_0[63]), .Z(n_19));
   OAI21_X1 i_84 (.A(n_196), .B1(n_195), .B2(n_21), .ZN(n_20));
   OAI21_X1 i_85 (.A(n_22), .B1(c[61]), .B2(p_0[61]), .ZN(n_21));
   NAND2_X1 i_86 (.A1(n_194), .A2(n_23), .ZN(n_22));
   AOI22_X1 i_87 (.A1(c[60]), .A2(p_0[60]), .B1(n_25), .B2(n_24), .ZN(n_23));
   XOR2_X1 i_88 (.A(c[60]), .B(p_0[60]), .Z(n_24));
   OAI21_X1 i_89 (.A(n_193), .B1(n_192), .B2(n_26), .ZN(n_25));
   OAI21_X1 i_90 (.A(n_27), .B1(c[58]), .B2(p_0[58]), .ZN(n_26));
   NAND2_X1 i_91 (.A1(n_191), .A2(n_28), .ZN(n_27));
   AOI22_X1 i_92 (.A1(c[57]), .A2(p_0[57]), .B1(n_189), .B2(n_29), .ZN(n_28));
   AOI21_X1 i_93 (.A(n_187), .B1(n_188), .B2(n_30), .ZN(n_29));
   AOI22_X1 i_94 (.A1(c[55]), .A2(p_0[55]), .B1(n_32), .B2(n_31), .ZN(n_30));
   XOR2_X1 i_95 (.A(c[55]), .B(p_0[55]), .Z(n_31));
   OAI21_X1 i_96 (.A(n_186), .B1(n_185), .B2(n_33), .ZN(n_32));
   OAI21_X1 i_97 (.A(n_34), .B1(c[53]), .B2(p_0[53]), .ZN(n_33));
   NAND2_X1 i_98 (.A1(n_184), .A2(n_35), .ZN(n_34));
   AOI22_X1 i_99 (.A1(c[52]), .A2(p_0[52]), .B1(n_182), .B2(n_36), .ZN(n_35));
   AOI21_X1 i_100 (.A(n_180), .B1(n_181), .B2(n_37), .ZN(n_36));
   AOI22_X1 i_101 (.A1(c[50]), .A2(p_0[50]), .B1(n_39), .B2(n_38), .ZN(n_37));
   XOR2_X1 i_102 (.A(c[50]), .B(p_0[50]), .Z(n_38));
   OAI21_X1 i_103 (.A(n_179), .B1(n_178), .B2(n_40), .ZN(n_39));
   OAI21_X1 i_104 (.A(n_41), .B1(c[48]), .B2(p_0[48]), .ZN(n_40));
   NAND2_X1 i_105 (.A1(n_177), .A2(n_42), .ZN(n_41));
   AOI22_X1 i_106 (.A1(c[47]), .A2(p_0[47]), .B1(n_175), .B2(n_43), .ZN(n_42));
   AOI21_X1 i_107 (.A(n_173), .B1(n_174), .B2(n_44), .ZN(n_43));
   AOI22_X1 i_108 (.A1(c[45]), .A2(p_0[45]), .B1(n_46), .B2(n_45), .ZN(n_44));
   XOR2_X1 i_109 (.A(c[45]), .B(p_0[45]), .Z(n_45));
   OAI21_X1 i_110 (.A(n_172), .B1(n_171), .B2(n_47), .ZN(n_46));
   OAI21_X1 i_111 (.A(n_48), .B1(c[43]), .B2(p_0[43]), .ZN(n_47));
   NAND2_X1 i_112 (.A1(n_170), .A2(n_49), .ZN(n_48));
   AOI22_X1 i_113 (.A1(c[42]), .A2(p_0[42]), .B1(n_168), .B2(n_50), .ZN(n_49));
   AOI21_X1 i_114 (.A(n_166), .B1(n_167), .B2(n_51), .ZN(n_50));
   AOI22_X1 i_115 (.A1(c[40]), .A2(p_0[40]), .B1(n_53), .B2(n_52), .ZN(n_51));
   XOR2_X1 i_116 (.A(c[40]), .B(p_0[40]), .Z(n_52));
   OAI21_X1 i_117 (.A(n_165), .B1(n_164), .B2(n_54), .ZN(n_53));
   OAI21_X1 i_118 (.A(n_55), .B1(c[38]), .B2(p_0[38]), .ZN(n_54));
   NAND2_X1 i_119 (.A1(n_163), .A2(n_56), .ZN(n_55));
   AOI22_X1 i_120 (.A1(c[37]), .A2(p_0[37]), .B1(n_161), .B2(n_57), .ZN(n_56));
   AOI21_X1 i_121 (.A(n_159), .B1(n_160), .B2(n_58), .ZN(n_57));
   AOI22_X1 i_122 (.A1(c[35]), .A2(p_0[35]), .B1(n_60), .B2(n_59), .ZN(n_58));
   XOR2_X1 i_123 (.A(c[35]), .B(p_0[35]), .Z(n_59));
   OAI21_X1 i_124 (.A(n_158), .B1(n_157), .B2(n_61), .ZN(n_60));
   OAI21_X1 i_125 (.A(n_62), .B1(c[33]), .B2(p_0[33]), .ZN(n_61));
   NAND2_X1 i_126 (.A1(n_156), .A2(n_63), .ZN(n_62));
   AOI22_X1 i_127 (.A1(c[32]), .A2(p_0[32]), .B1(n_154), .B2(n_64), .ZN(n_63));
   AOI21_X1 i_128 (.A(n_152), .B1(n_153), .B2(n_65), .ZN(n_64));
   AOI22_X1 i_129 (.A1(c[30]), .A2(p_0[30]), .B1(n_67), .B2(n_66), .ZN(n_65));
   XOR2_X1 i_130 (.A(c[30]), .B(p_0[30]), .Z(n_66));
   OAI21_X1 i_131 (.A(n_151), .B1(n_150), .B2(n_68), .ZN(n_67));
   OAI21_X1 i_132 (.A(n_69), .B1(c[28]), .B2(p_0[28]), .ZN(n_68));
   NAND2_X1 i_133 (.A1(n_149), .A2(n_70), .ZN(n_69));
   AOI22_X1 i_134 (.A1(c[27]), .A2(p_0[27]), .B1(n_147), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_135 (.A(n_145), .B1(n_146), .B2(n_72), .ZN(n_71));
   AOI22_X1 i_136 (.A1(c[25]), .A2(p_0[25]), .B1(n_74), .B2(n_73), .ZN(n_72));
   XOR2_X1 i_137 (.A(c[25]), .B(p_0[25]), .Z(n_73));
   OAI21_X1 i_138 (.A(n_144), .B1(n_143), .B2(n_75), .ZN(n_74));
   OAI21_X1 i_139 (.A(n_76), .B1(c[23]), .B2(p_0[23]), .ZN(n_75));
   NAND2_X1 i_140 (.A1(n_142), .A2(n_77), .ZN(n_76));
   AOI22_X1 i_141 (.A1(c[22]), .A2(p_0[22]), .B1(n_140), .B2(n_78), .ZN(n_77));
   AOI21_X1 i_142 (.A(n_138), .B1(n_139), .B2(n_79), .ZN(n_78));
   AOI22_X1 i_143 (.A1(c[20]), .A2(p_0[20]), .B1(n_81), .B2(n_80), .ZN(n_79));
   XOR2_X1 i_144 (.A(c[20]), .B(p_0[20]), .Z(n_80));
   INV_X1 i_145 (.A(n_82), .ZN(n_81));
   AOI22_X1 i_146 (.A1(c[19]), .A2(p_0[19]), .B1(n_84), .B2(n_83), .ZN(n_82));
   XOR2_X1 i_147 (.A(c[19]), .B(p_0[19]), .Z(n_83));
   INV_X1 i_148 (.A(n_85), .ZN(n_84));
   AOI22_X1 i_149 (.A1(c[18]), .A2(p_0[18]), .B1(n_87), .B2(n_86), .ZN(n_85));
   XOR2_X1 i_150 (.A(c[18]), .B(p_0[18]), .Z(n_86));
   INV_X1 i_151 (.A(n_88), .ZN(n_87));
   AOI22_X1 i_152 (.A1(c[17]), .A2(p_0[17]), .B1(n_136), .B2(n_89), .ZN(n_88));
   OAI21_X1 i_153 (.A(n_90), .B1(n_202), .B2(n_199), .ZN(n_89));
   OAI21_X1 i_154 (.A(n_91), .B1(c[16]), .B2(p_0[16]), .ZN(n_90));
   OAI21_X1 i_155 (.A(n_135), .B1(n_93), .B2(n_92), .ZN(n_91));
   OAI21_X1 i_156 (.A(n_135), .B1(c[15]), .B2(p_0[15]), .ZN(n_92));
   AOI22_X1 i_157 (.A1(c[14]), .A2(p_0[14]), .B1(n_95), .B2(n_94), .ZN(n_93));
   XOR2_X1 i_158 (.A(c[14]), .B(p_0[14]), .Z(n_94));
   INV_X1 i_159 (.A(n_96), .ZN(n_95));
   AOI22_X1 i_160 (.A1(c[13]), .A2(p_0[13]), .B1(n_98), .B2(n_97), .ZN(n_96));
   XOR2_X1 i_161 (.A(c[13]), .B(p_0[13]), .Z(n_97));
   INV_X1 i_162 (.A(n_99), .ZN(n_98));
   AOI22_X1 i_163 (.A1(c[12]), .A2(p_0[12]), .B1(n_101), .B2(n_100), .ZN(n_99));
   XOR2_X1 i_164 (.A(c[12]), .B(p_0[12]), .Z(n_100));
   INV_X1 i_165 (.A(n_102), .ZN(n_101));
   AOI22_X1 i_166 (.A1(c[11]), .A2(p_0[11]), .B1(n_104), .B2(n_103), .ZN(n_102));
   XOR2_X1 i_167 (.A(c[11]), .B(p_0[11]), .Z(n_103));
   INV_X1 i_168 (.A(n_105), .ZN(n_104));
   AOI22_X1 i_169 (.A1(c[10]), .A2(p_0[10]), .B1(n_107), .B2(n_106), .ZN(n_105));
   XOR2_X1 i_170 (.A(c[10]), .B(p_0[10]), .Z(n_106));
   INV_X1 i_171 (.A(n_108), .ZN(n_107));
   AOI22_X1 i_172 (.A1(c[9]), .A2(p_0[9]), .B1(n_110), .B2(n_109), .ZN(n_108));
   XOR2_X1 i_173 (.A(c[9]), .B(p_0[9]), .Z(n_109));
   INV_X1 i_174 (.A(n_111), .ZN(n_110));
   AOI22_X1 i_175 (.A1(c[8]), .A2(p_0[8]), .B1(n_113), .B2(n_112), .ZN(n_111));
   XOR2_X1 i_176 (.A(c[8]), .B(p_0[8]), .Z(n_112));
   INV_X1 i_177 (.A(n_114), .ZN(n_113));
   AOI22_X1 i_178 (.A1(c[7]), .A2(p_0[7]), .B1(n_116), .B2(n_115), .ZN(n_114));
   XOR2_X1 i_179 (.A(c[7]), .B(p_0[7]), .Z(n_115));
   INV_X1 i_180 (.A(n_117), .ZN(n_116));
   AOI22_X1 i_181 (.A1(c[6]), .A2(p_0[6]), .B1(n_119), .B2(n_118), .ZN(n_117));
   XOR2_X1 i_182 (.A(c[6]), .B(p_0[6]), .Z(n_118));
   INV_X1 i_183 (.A(n_120), .ZN(n_119));
   AOI22_X1 i_184 (.A1(c[5]), .A2(p_0[5]), .B1(n_122), .B2(n_121), .ZN(n_120));
   XOR2_X1 i_185 (.A(c[5]), .B(p_0[5]), .Z(n_121));
   INV_X1 i_186 (.A(n_123), .ZN(n_122));
   AOI22_X1 i_187 (.A1(c[4]), .A2(p_0[4]), .B1(n_125), .B2(n_124), .ZN(n_123));
   XOR2_X1 i_188 (.A(c[4]), .B(p_0[4]), .Z(n_124));
   INV_X1 i_189 (.A(n_126), .ZN(n_125));
   AOI22_X1 i_190 (.A1(c[3]), .A2(p_0[3]), .B1(n_128), .B2(n_127), .ZN(n_126));
   XOR2_X1 i_191 (.A(c[3]), .B(p_0[3]), .Z(n_127));
   INV_X1 i_192 (.A(n_129), .ZN(n_128));
   AOI22_X1 i_193 (.A1(c[2]), .A2(p_0[2]), .B1(n_133), .B2(n_130), .ZN(n_129));
   AOI21_X1 i_194 (.A(n_131), .B1(n_201), .B2(n_198), .ZN(n_130));
   AOI21_X1 i_195 (.A(n_132), .B1(c[1]), .B2(p_0[1]), .ZN(n_131));
   NOR2_X1 i_196 (.A1(n_200), .A2(n_197), .ZN(n_132));
   INV_X1 i_197 (.A(n_134), .ZN(n_133));
   XNOR2_X1 i_198 (.A(c[2]), .B(p_0[2]), .ZN(n_134));
   NAND2_X1 i_199 (.A1(c[15]), .A2(p_0[15]), .ZN(n_135));
   INV_X1 i_200 (.A(n_137), .ZN(n_136));
   XNOR2_X1 i_201 (.A(c[17]), .B(p_0[17]), .ZN(n_137));
   NOR2_X1 i_202 (.A1(c[21]), .A2(p_0[21]), .ZN(n_138));
   NAND2_X1 i_203 (.A1(c[21]), .A2(p_0[21]), .ZN(n_139));
   INV_X1 i_204 (.A(n_141), .ZN(n_140));
   XNOR2_X1 i_205 (.A(c[22]), .B(p_0[22]), .ZN(n_141));
   NAND2_X1 i_206 (.A1(c[23]), .A2(p_0[23]), .ZN(n_142));
   OAI21_X1 i_207 (.A(n_144), .B1(c[24]), .B2(p_0[24]), .ZN(n_143));
   NAND2_X1 i_208 (.A1(c[24]), .A2(p_0[24]), .ZN(n_144));
   NOR2_X1 i_209 (.A1(c[26]), .A2(p_0[26]), .ZN(n_145));
   NAND2_X1 i_210 (.A1(c[26]), .A2(p_0[26]), .ZN(n_146));
   INV_X1 i_211 (.A(n_148), .ZN(n_147));
   XNOR2_X1 i_212 (.A(c[27]), .B(p_0[27]), .ZN(n_148));
   NAND2_X1 i_213 (.A1(c[28]), .A2(p_0[28]), .ZN(n_149));
   OAI21_X1 i_214 (.A(n_151), .B1(c[29]), .B2(p_0[29]), .ZN(n_150));
   NAND2_X1 i_215 (.A1(c[29]), .A2(p_0[29]), .ZN(n_151));
   NOR2_X1 i_216 (.A1(c[31]), .A2(p_0[31]), .ZN(n_152));
   NAND2_X1 i_217 (.A1(c[31]), .A2(p_0[31]), .ZN(n_153));
   INV_X1 i_218 (.A(n_155), .ZN(n_154));
   XNOR2_X1 i_219 (.A(c[32]), .B(p_0[32]), .ZN(n_155));
   NAND2_X1 i_220 (.A1(c[33]), .A2(p_0[33]), .ZN(n_156));
   OAI21_X1 i_221 (.A(n_158), .B1(c[34]), .B2(p_0[34]), .ZN(n_157));
   NAND2_X1 i_222 (.A1(c[34]), .A2(p_0[34]), .ZN(n_158));
   NOR2_X1 i_223 (.A1(c[36]), .A2(p_0[36]), .ZN(n_159));
   NAND2_X1 i_224 (.A1(c[36]), .A2(p_0[36]), .ZN(n_160));
   INV_X1 i_225 (.A(n_162), .ZN(n_161));
   XNOR2_X1 i_226 (.A(c[37]), .B(p_0[37]), .ZN(n_162));
   NAND2_X1 i_227 (.A1(c[38]), .A2(p_0[38]), .ZN(n_163));
   OAI21_X1 i_228 (.A(n_165), .B1(c[39]), .B2(p_0[39]), .ZN(n_164));
   NAND2_X1 i_229 (.A1(c[39]), .A2(p_0[39]), .ZN(n_165));
   NOR2_X1 i_230 (.A1(c[41]), .A2(p_0[41]), .ZN(n_166));
   NAND2_X1 i_231 (.A1(c[41]), .A2(p_0[41]), .ZN(n_167));
   INV_X1 i_232 (.A(n_169), .ZN(n_168));
   XNOR2_X1 i_233 (.A(c[42]), .B(p_0[42]), .ZN(n_169));
   NAND2_X1 i_234 (.A1(c[43]), .A2(p_0[43]), .ZN(n_170));
   OAI21_X1 i_235 (.A(n_172), .B1(c[44]), .B2(p_0[44]), .ZN(n_171));
   NAND2_X1 i_236 (.A1(c[44]), .A2(p_0[44]), .ZN(n_172));
   NOR2_X1 i_237 (.A1(c[46]), .A2(p_0[46]), .ZN(n_173));
   NAND2_X1 i_238 (.A1(c[46]), .A2(p_0[46]), .ZN(n_174));
   INV_X1 i_239 (.A(n_176), .ZN(n_175));
   XNOR2_X1 i_240 (.A(c[47]), .B(p_0[47]), .ZN(n_176));
   NAND2_X1 i_241 (.A1(c[48]), .A2(p_0[48]), .ZN(n_177));
   OAI21_X1 i_242 (.A(n_179), .B1(c[49]), .B2(p_0[49]), .ZN(n_178));
   NAND2_X1 i_243 (.A1(c[49]), .A2(p_0[49]), .ZN(n_179));
   NOR2_X1 i_244 (.A1(c[51]), .A2(p_0[51]), .ZN(n_180));
   NAND2_X1 i_245 (.A1(c[51]), .A2(p_0[51]), .ZN(n_181));
   INV_X1 i_246 (.A(n_183), .ZN(n_182));
   XNOR2_X1 i_247 (.A(c[52]), .B(p_0[52]), .ZN(n_183));
   NAND2_X1 i_248 (.A1(c[53]), .A2(p_0[53]), .ZN(n_184));
   OAI21_X1 i_249 (.A(n_186), .B1(c[54]), .B2(p_0[54]), .ZN(n_185));
   NAND2_X1 i_250 (.A1(c[54]), .A2(p_0[54]), .ZN(n_186));
   NOR2_X1 i_251 (.A1(c[56]), .A2(p_0[56]), .ZN(n_187));
   NAND2_X1 i_252 (.A1(c[56]), .A2(p_0[56]), .ZN(n_188));
   INV_X1 i_253 (.A(n_190), .ZN(n_189));
   XNOR2_X1 i_254 (.A(c[57]), .B(p_0[57]), .ZN(n_190));
   NAND2_X1 i_255 (.A1(c[58]), .A2(p_0[58]), .ZN(n_191));
   OAI21_X1 i_256 (.A(n_193), .B1(c[59]), .B2(p_0[59]), .ZN(n_192));
   NAND2_X1 i_257 (.A1(c[59]), .A2(p_0[59]), .ZN(n_193));
   NAND2_X1 i_258 (.A1(c[61]), .A2(p_0[61]), .ZN(n_194));
   OAI21_X1 i_259 (.A(n_196), .B1(c[62]), .B2(p_0[62]), .ZN(n_195));
   NAND2_X1 i_260 (.A1(c[62]), .A2(p_0[62]), .ZN(n_196));
   INV_X1 i_261 (.A(p_0[0]), .ZN(n_197));
   INV_X1 i_262 (.A(p_0[1]), .ZN(n_198));
   INV_X1 i_263 (.A(p_0[16]), .ZN(n_199));
   INV_X1 i_264 (.A(c[0]), .ZN(n_200));
   INV_X1 i_265 (.A(c[1]), .ZN(n_201));
   INV_X1 i_266 (.A(c[16]), .ZN(n_202));
endmodule

module Radix4(a, b, read_data3, clk, start, start_shift, start_i);
   input [31:0]a;
   input [31:0]b;
   output [63:0]read_data3;
   input clk;
   input start;
   input [4:0]start_shift;
   input [4:0]start_i;

   wire [31:0]read_data2;
   wire [31:0]read_data;
   wire n_0_0;
   wire [63:0]res;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_1;
   wire n_0_0_2;
   wire n_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_3;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_66;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_67;
   wire n_0_0_17;
   wire n_0_68;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_70;
   wire n_0_0_20;
   wire n_0_71;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_72;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_73;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_74;
   wire n_0_0_33;
   wire n_0_75;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_105;
   wire n_0_0_38;
   wire n_0_69;
   wire n_0_0_39;
   wire n_0_235;
   wire n_0_0_40;
   wire n_0_236;
   wire n_0_0_41;
   wire n_0_237;
   wire n_0_0_42;
   wire n_0_238;
   wire n_0_0_43;
   wire n_0_239;
   wire n_0_0_44;
   wire n_0_240;
   wire n_0_0_45;
   wire n_0_241;
   wire n_0_0_46;
   wire n_0_242;
   wire n_0_0_47;
   wire n_0_243;
   wire n_0_0_48;
   wire n_0_244;
   wire n_0_0_49;
   wire n_0_245;
   wire n_0_0_50;
   wire n_0_246;
   wire n_0_0_51;
   wire n_0_247;
   wire n_0_0_52;
   wire n_0_248;
   wire n_0_0_53;
   wire n_0_249;
   wire n_0_0_54;
   wire n_0_250;
   wire n_0_0_55;
   wire n_0_251;
   wire n_0_0_56;
   wire n_0_252;
   wire n_0_0_57;
   wire n_0_253;
   wire n_0_0_58;
   wire n_0_254;
   wire n_0_0_59;
   wire n_0_255;
   wire n_0_0_60;
   wire n_0_256;
   wire n_0_0_61;
   wire n_0_257;
   wire n_0_0_62;
   wire n_0_258;
   wire n_0_0_63;
   wire n_0_259;
   wire n_0_0_64;
   wire n_0_260;
   wire n_0_0_65;
   wire n_0_261;
   wire n_0_0_66;
   wire n_0_262;
   wire n_0_0_67;
   wire n_0_263;
   wire n_0_0_68;
   wire n_0_264;
   wire n_0_0_69;
   wire n_0_265;
   wire n_0_0_70;
   wire n_0_266;
   wire n_0_0_71;
   wire n_0_267;
   wire n_0_0_72;
   wire n_0_268;
   wire n_0_0_73;
   wire n_0_269;
   wire n_0_0_74;
   wire n_0_76;
   wire n_0_0_75;
   wire n_0_77;
   wire n_0_0_76;
   wire n_0_78;
   wire n_0_0_77;
   wire n_0_79;
   wire n_0_0_78;
   wire n_0_80;
   wire n_0_0_79;
   wire n_0_81;
   wire n_0_0_80;
   wire n_0_82;
   wire n_0_0_81;
   wire n_0_83;
   wire n_0_0_82;
   wire n_0_84;
   wire n_0_0_83;
   wire n_0_85;
   wire n_0_0_84;
   wire n_0_86;
   wire n_0_0_85;
   wire n_0_87;
   wire n_0_0_86;
   wire n_0_88;
   wire n_0_0_87;
   wire n_0_89;
   wire n_0_0_88;
   wire n_0_90;
   wire n_0_0_89;
   wire n_0_91;
   wire n_0_0_90;
   wire n_0_92;
   wire n_0_0_91;
   wire n_0_93;
   wire n_0_0_92;
   wire n_0_94;
   wire n_0_0_93;
   wire n_0_95;
   wire n_0_0_94;
   wire n_0_96;
   wire n_0_0_95;
   wire n_0_97;
   wire n_0_0_96;
   wire n_0_98;
   wire n_0_0_97;
   wire n_0_99;
   wire n_0_0_98;
   wire n_0_100;
   wire n_0_0_99;
   wire n_0_101;
   wire n_0_0_100;
   wire n_0_102;
   wire n_0_0_101;
   wire n_0_103;
   wire n_0_0_102;
   wire n_0_104;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_108;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_109;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_110;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_111;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_112;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_113;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_114;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_115;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_116;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_117;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_118;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_119;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_120;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_121;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_122;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_123;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_124;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_125;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_126;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_127;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_128;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_129;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_130;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_131;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_132;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_133;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_134;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_135;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_136;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_137;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_138;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_139;
   wire n_0_0_422;
   wire n_0_107;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_140;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_141;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_142;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_143;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_144;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_145;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_146;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_147;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_148;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_149;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_150;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_151;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_152;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_153;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_154;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_155;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_156;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_157;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_158;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_159;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_160;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_161;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_162;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_163;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_164;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_165;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_166;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_167;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_168;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_169;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_170;
   wire write_en;
   wire [63:0]c;
   wire [5:0]shift;
   wire [5:0]i;
   wire n_0_106;

   regFile r (.read_data(read_data), .read_data2(read_data2), .write_en(write_en), 
      .write_data(a), .write_data2(b), .clk(clk));
   regFile64 r2 (.read_data(read_data3), .write_en(), .write_data(res), .clk(clk));
   CLKGATETST_X1 clk_gate_res_reg (.CK(clk), .E(n_0_105), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \res_reg[63]  (.D(n_0_234), .CK(n_0_0), .Q(res[63]), .QN());
   DFF_X1 \res_reg[62]  (.D(n_0_233), .CK(n_0_0), .Q(res[62]), .QN());
   DFF_X1 \res_reg[61]  (.D(n_0_232), .CK(n_0_0), .Q(res[61]), .QN());
   DFF_X1 \res_reg[60]  (.D(n_0_231), .CK(n_0_0), .Q(res[60]), .QN());
   DFF_X1 \res_reg[59]  (.D(n_0_230), .CK(n_0_0), .Q(res[59]), .QN());
   DFF_X1 \res_reg[58]  (.D(n_0_229), .CK(n_0_0), .Q(res[58]), .QN());
   DFF_X1 \res_reg[57]  (.D(n_0_228), .CK(n_0_0), .Q(res[57]), .QN());
   DFF_X1 \res_reg[56]  (.D(n_0_227), .CK(n_0_0), .Q(res[56]), .QN());
   DFF_X1 \res_reg[55]  (.D(n_0_226), .CK(n_0_0), .Q(res[55]), .QN());
   DFF_X1 \res_reg[54]  (.D(n_0_225), .CK(n_0_0), .Q(res[54]), .QN());
   DFF_X1 \res_reg[53]  (.D(n_0_224), .CK(n_0_0), .Q(res[53]), .QN());
   DFF_X1 \res_reg[52]  (.D(n_0_223), .CK(n_0_0), .Q(res[52]), .QN());
   DFF_X1 \res_reg[51]  (.D(n_0_222), .CK(n_0_0), .Q(res[51]), .QN());
   DFF_X1 \res_reg[50]  (.D(n_0_221), .CK(n_0_0), .Q(res[50]), .QN());
   DFF_X1 \res_reg[49]  (.D(n_0_220), .CK(n_0_0), .Q(res[49]), .QN());
   DFF_X1 \res_reg[48]  (.D(n_0_219), .CK(n_0_0), .Q(res[48]), .QN());
   DFF_X1 \res_reg[47]  (.D(n_0_218), .CK(n_0_0), .Q(res[47]), .QN());
   DFF_X1 \res_reg[46]  (.D(n_0_217), .CK(n_0_0), .Q(res[46]), .QN());
   DFF_X1 \res_reg[45]  (.D(n_0_216), .CK(n_0_0), .Q(res[45]), .QN());
   DFF_X1 \res_reg[44]  (.D(n_0_215), .CK(n_0_0), .Q(res[44]), .QN());
   DFF_X1 \res_reg[43]  (.D(n_0_214), .CK(n_0_0), .Q(res[43]), .QN());
   DFF_X1 \res_reg[42]  (.D(n_0_213), .CK(n_0_0), .Q(res[42]), .QN());
   DFF_X1 \res_reg[41]  (.D(n_0_212), .CK(n_0_0), .Q(res[41]), .QN());
   DFF_X1 \res_reg[40]  (.D(n_0_211), .CK(n_0_0), .Q(res[40]), .QN());
   DFF_X1 \res_reg[39]  (.D(n_0_210), .CK(n_0_0), .Q(res[39]), .QN());
   DFF_X1 \res_reg[38]  (.D(n_0_209), .CK(n_0_0), .Q(res[38]), .QN());
   DFF_X1 \res_reg[37]  (.D(n_0_208), .CK(n_0_0), .Q(res[37]), .QN());
   DFF_X1 \res_reg[36]  (.D(n_0_207), .CK(n_0_0), .Q(res[36]), .QN());
   DFF_X1 \res_reg[35]  (.D(n_0_206), .CK(n_0_0), .Q(res[35]), .QN());
   DFF_X1 \res_reg[34]  (.D(n_0_205), .CK(n_0_0), .Q(res[34]), .QN());
   DFF_X1 \res_reg[33]  (.D(n_0_204), .CK(n_0_0), .Q(res[33]), .QN());
   DFF_X1 \res_reg[32]  (.D(n_0_203), .CK(n_0_0), .Q(res[32]), .QN());
   DFF_X1 \res_reg[31]  (.D(n_0_202), .CK(n_0_0), .Q(res[31]), .QN());
   DFF_X1 \res_reg[30]  (.D(n_0_201), .CK(n_0_0), .Q(res[30]), .QN());
   DFF_X1 \res_reg[29]  (.D(n_0_200), .CK(n_0_0), .Q(res[29]), .QN());
   DFF_X1 \res_reg[28]  (.D(n_0_199), .CK(n_0_0), .Q(res[28]), .QN());
   DFF_X1 \res_reg[27]  (.D(n_0_198), .CK(n_0_0), .Q(res[27]), .QN());
   DFF_X1 \res_reg[26]  (.D(n_0_197), .CK(n_0_0), .Q(res[26]), .QN());
   DFF_X1 \res_reg[25]  (.D(n_0_196), .CK(n_0_0), .Q(res[25]), .QN());
   DFF_X1 \res_reg[24]  (.D(n_0_195), .CK(n_0_0), .Q(res[24]), .QN());
   DFF_X1 \res_reg[23]  (.D(n_0_194), .CK(n_0_0), .Q(res[23]), .QN());
   DFF_X1 \res_reg[22]  (.D(n_0_193), .CK(n_0_0), .Q(res[22]), .QN());
   DFF_X1 \res_reg[21]  (.D(n_0_192), .CK(n_0_0), .Q(res[21]), .QN());
   DFF_X1 \res_reg[20]  (.D(n_0_191), .CK(n_0_0), .Q(res[20]), .QN());
   DFF_X1 \res_reg[19]  (.D(n_0_190), .CK(n_0_0), .Q(res[19]), .QN());
   DFF_X1 \res_reg[18]  (.D(n_0_189), .CK(n_0_0), .Q(res[18]), .QN());
   DFF_X1 \res_reg[17]  (.D(n_0_188), .CK(n_0_0), .Q(res[17]), .QN());
   DFF_X1 \res_reg[16]  (.D(n_0_187), .CK(n_0_0), .Q(res[16]), .QN());
   DFF_X1 \res_reg[15]  (.D(n_0_186), .CK(n_0_0), .Q(res[15]), .QN());
   DFF_X1 \res_reg[14]  (.D(n_0_185), .CK(n_0_0), .Q(res[14]), .QN());
   DFF_X1 \res_reg[13]  (.D(n_0_184), .CK(n_0_0), .Q(res[13]), .QN());
   DFF_X1 \res_reg[12]  (.D(n_0_183), .CK(n_0_0), .Q(res[12]), .QN());
   DFF_X1 \res_reg[11]  (.D(n_0_182), .CK(n_0_0), .Q(res[11]), .QN());
   DFF_X1 \res_reg[10]  (.D(n_0_181), .CK(n_0_0), .Q(res[10]), .QN());
   DFF_X1 \res_reg[9]  (.D(n_0_180), .CK(n_0_0), .Q(res[9]), .QN());
   DFF_X1 \res_reg[8]  (.D(n_0_179), .CK(n_0_0), .Q(res[8]), .QN());
   DFF_X1 \res_reg[7]  (.D(n_0_178), .CK(n_0_0), .Q(res[7]), .QN());
   DFF_X1 \res_reg[6]  (.D(n_0_177), .CK(n_0_0), .Q(res[6]), .QN());
   DFF_X1 \res_reg[5]  (.D(n_0_176), .CK(n_0_0), .Q(res[5]), .QN());
   DFF_X1 \res_reg[4]  (.D(n_0_175), .CK(n_0_0), .Q(res[4]), .QN());
   DFF_X1 \res_reg[3]  (.D(n_0_174), .CK(n_0_0), .Q(res[3]), .QN());
   DFF_X1 \res_reg[2]  (.D(n_0_173), .CK(n_0_0), .Q(res[2]), .QN());
   DFF_X1 \res_reg[1]  (.D(n_0_172), .CK(n_0_0), .Q(res[1]), .QN());
   DFF_X1 \res_reg[0]  (.D(n_0_171), .CK(n_0_0), .Q(res[0]), .QN());
   datapath i_0_3 (.p_0({n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
      n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, uc_0}), .read_data2(read_data2));
   datapath__0_128 i_0_4 (.p_0({uc_1, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, 
      n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, 
      n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, 
      n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, uc_2}), 
      .p_1({1'b0, read_data2[31], read_data2[30], read_data2[29], read_data2[28], 
      read_data2[27], read_data2[26], read_data2[25], read_data2[24], 
      read_data2[23], read_data2[22], read_data2[21], read_data2[20], 
      read_data2[19], read_data2[18], read_data2[17], read_data2[16], 
      read_data2[15], read_data2[14], read_data2[13], read_data2[12], 
      read_data2[11], read_data2[10], read_data2[9], read_data2[8], 
      read_data2[7], read_data2[6], read_data2[5], read_data2[4], read_data2[3], 
      read_data2[2], read_data2[1], read_data2[0]}));
   datapath__0_142 i_0_11 (.c(c), .p_0({n_0_107, n_0_170, n_0_169, n_0_168, 
      n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, 
      n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, 
      n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, 
      n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, 
      n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, 
      n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108}), .p_1({n_0_234, n_0_233, n_0_232, 
      n_0_231, n_0_230, n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, 
      n_0_223, n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, 
      n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, 
      n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, 
      n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, n_0_192, 
      n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, 
      n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, 
      n_0_175, n_0_174, n_0_173, n_0_172, n_0_171}));
   NAND2_X1 i_0_0_0 (.A1(start_i[0]), .A2(start), .ZN(n_0_0_0));
   INV_X1 i_0_0_1 (.A(i[0]), .ZN(n_0_0_1));
   OAI21_X1 i_0_0_2 (.A(n_0_0_0), .B1(n_0_0_1), .B2(start), .ZN(n_0_1));
   NAND2_X1 i_0_0_3 (.A1(start_i[1]), .A2(start), .ZN(n_0_0_2));
   OAI21_X1 i_0_0_4 (.A(n_0_0_2), .B1(start), .B2(i[1]), .ZN(n_0_2));
   NAND2_X1 i_0_0_5 (.A1(start_i[2]), .A2(start), .ZN(n_0_0_3));
   INV_X1 i_0_0_6 (.A(start), .ZN(n_0_0_4));
   OAI21_X1 i_0_0_7 (.A(n_0_0_4), .B1(i[1]), .B2(i[2]), .ZN(n_0_0_5));
   INV_X1 i_0_0_8 (.A(i[1]), .ZN(n_0_0_6));
   INV_X1 i_0_0_9 (.A(i[2]), .ZN(n_0_0_7));
   NOR2_X1 i_0_0_10 (.A1(n_0_0_6), .A2(n_0_0_7), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_11 (.A(n_0_0_3), .B1(n_0_0_5), .B2(n_0_0_8), .ZN(n_0_3));
   NAND2_X1 i_0_0_12 (.A1(n_0_0_8), .A2(i[3]), .ZN(n_0_0_9));
   OAI21_X1 i_0_0_13 (.A(n_0_0_9), .B1(i[3]), .B2(n_0_0_8), .ZN(n_0_0_10));
   INV_X1 i_0_0_14 (.A(start_i[3]), .ZN(n_0_0_11));
   AOI22_X1 i_0_0_15 (.A1(n_0_0_10), .A2(n_0_0_4), .B1(n_0_0_11), .B2(start), 
      .ZN(n_0_66));
   NAND2_X1 i_0_0_16 (.A1(start_i[4]), .A2(start), .ZN(n_0_0_12));
   INV_X1 i_0_0_17 (.A(n_0_0_9), .ZN(n_0_0_13));
   OAI21_X1 i_0_0_18 (.A(n_0_0_4), .B1(n_0_0_13), .B2(i[4]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_19 (.A1(n_0_0_13), .A2(i[4]), .ZN(n_0_0_15));
   INV_X1 i_0_0_20 (.A(n_0_0_15), .ZN(n_0_0_16));
   OAI21_X1 i_0_0_21 (.A(n_0_0_12), .B1(n_0_0_14), .B2(n_0_0_16), .ZN(n_0_67));
   INV_X1 i_0_0_22 (.A(i[5]), .ZN(n_0_0_17));
   AOI221_X1 i_0_0_23 (.A(start), .B1(n_0_0_16), .B2(i[5]), .C1(n_0_0_17), 
      .C2(n_0_0_15), .ZN(n_0_68));
   NAND2_X1 i_0_0_24 (.A1(start_shift[0]), .A2(start), .ZN(n_0_0_18));
   INV_X1 i_0_0_25 (.A(shift[0]), .ZN(n_0_0_19));
   OAI21_X1 i_0_0_26 (.A(n_0_0_18), .B1(n_0_0_19), .B2(start), .ZN(n_0_70));
   NAND2_X1 i_0_0_27 (.A1(start_shift[1]), .A2(start), .ZN(n_0_0_20));
   OAI21_X1 i_0_0_28 (.A(n_0_0_20), .B1(start), .B2(shift[1]), .ZN(n_0_71));
   NAND2_X1 i_0_0_29 (.A1(start_shift[2]), .A2(start), .ZN(n_0_0_21));
   OAI21_X1 i_0_0_30 (.A(n_0_0_4), .B1(shift[2]), .B2(shift[1]), .ZN(n_0_0_22));
   INV_X1 i_0_0_31 (.A(shift[2]), .ZN(n_0_0_23));
   INV_X1 i_0_0_32 (.A(shift[1]), .ZN(n_0_0_24));
   NOR2_X1 i_0_0_33 (.A1(n_0_0_23), .A2(n_0_0_24), .ZN(n_0_0_25));
   OAI21_X1 i_0_0_34 (.A(n_0_0_21), .B1(n_0_0_22), .B2(n_0_0_25), .ZN(n_0_72));
   NAND2_X1 i_0_0_35 (.A1(start_shift[3]), .A2(start), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_36 (.A(n_0_0_4), .B1(n_0_0_25), .B2(shift[3]), .ZN(n_0_0_27));
   AND2_X1 i_0_0_37 (.A1(n_0_0_25), .A2(shift[3]), .ZN(n_0_0_28));
   OAI21_X1 i_0_0_38 (.A(n_0_0_26), .B1(n_0_0_27), .B2(n_0_0_28), .ZN(n_0_73));
   NAND2_X1 i_0_0_39 (.A1(start_shift[4]), .A2(start), .ZN(n_0_0_29));
   OAI21_X1 i_0_0_40 (.A(n_0_0_4), .B1(n_0_0_28), .B2(shift[4]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_28), .A2(shift[4]), .ZN(n_0_0_31));
   INV_X1 i_0_0_42 (.A(n_0_0_31), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_43 (.A(n_0_0_29), .B1(n_0_0_30), .B2(n_0_0_32), .ZN(n_0_74));
   INV_X1 i_0_0_44 (.A(shift[5]), .ZN(n_0_0_33));
   AOI221_X1 i_0_0_45 (.A(start), .B1(n_0_0_32), .B2(shift[5]), .C1(n_0_0_33), 
      .C2(n_0_0_31), .ZN(n_0_75));
   NOR2_X1 i_0_0_46 (.A1(i[0]), .A2(i[2]), .ZN(n_0_0_34));
   NOR2_X1 i_0_0_47 (.A1(i[4]), .A2(i[3]), .ZN(n_0_0_35));
   NAND3_X1 i_0_0_48 (.A1(n_0_0_34), .A2(n_0_0_35), .A3(n_0_0_6), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_49 (.A1(n_0_0_36), .A2(i[5]), .ZN(n_0_0_37));
   AND2_X1 i_0_0_50 (.A1(n_0_0_37), .A2(n_0_0_4), .ZN(n_0_105));
   NOR2_X1 i_0_0_51 (.A1(n_0_0_37), .A2(start), .ZN(n_0_0_38));
   INV_X1 i_0_0_52 (.A(n_0_0_38), .ZN(n_0_69));
   AOI22_X1 i_0_0_53 (.A1(n_0_105), .A2(n_0_171), .B1(n_0_0_38), .B2(res[0]), 
      .ZN(n_0_0_39));
   INV_X1 i_0_0_54 (.A(n_0_0_39), .ZN(n_0_235));
   AOI22_X1 i_0_0_55 (.A1(n_0_105), .A2(n_0_172), .B1(n_0_0_38), .B2(res[1]), 
      .ZN(n_0_0_40));
   INV_X1 i_0_0_56 (.A(n_0_0_40), .ZN(n_0_236));
   AOI22_X1 i_0_0_57 (.A1(n_0_105), .A2(n_0_173), .B1(n_0_0_38), .B2(res[2]), 
      .ZN(n_0_0_41));
   INV_X1 i_0_0_58 (.A(n_0_0_41), .ZN(n_0_237));
   AOI22_X1 i_0_0_59 (.A1(n_0_105), .A2(n_0_174), .B1(n_0_0_38), .B2(res[3]), 
      .ZN(n_0_0_42));
   INV_X1 i_0_0_60 (.A(n_0_0_42), .ZN(n_0_238));
   AOI22_X1 i_0_0_61 (.A1(n_0_105), .A2(n_0_175), .B1(n_0_0_38), .B2(res[4]), 
      .ZN(n_0_0_43));
   INV_X1 i_0_0_62 (.A(n_0_0_43), .ZN(n_0_239));
   AOI22_X1 i_0_0_63 (.A1(n_0_105), .A2(n_0_176), .B1(n_0_0_38), .B2(res[5]), 
      .ZN(n_0_0_44));
   INV_X1 i_0_0_64 (.A(n_0_0_44), .ZN(n_0_240));
   AOI22_X1 i_0_0_65 (.A1(n_0_105), .A2(n_0_177), .B1(n_0_0_38), .B2(res[6]), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_66 (.A(n_0_0_45), .ZN(n_0_241));
   AOI22_X1 i_0_0_67 (.A1(n_0_105), .A2(n_0_178), .B1(n_0_0_38), .B2(res[7]), 
      .ZN(n_0_0_46));
   INV_X1 i_0_0_68 (.A(n_0_0_46), .ZN(n_0_242));
   AOI22_X1 i_0_0_69 (.A1(n_0_105), .A2(n_0_179), .B1(n_0_0_38), .B2(res[8]), 
      .ZN(n_0_0_47));
   INV_X1 i_0_0_70 (.A(n_0_0_47), .ZN(n_0_243));
   AOI22_X1 i_0_0_71 (.A1(n_0_105), .A2(n_0_180), .B1(n_0_0_38), .B2(res[9]), 
      .ZN(n_0_0_48));
   INV_X1 i_0_0_72 (.A(n_0_0_48), .ZN(n_0_244));
   AOI22_X1 i_0_0_73 (.A1(n_0_105), .A2(n_0_181), .B1(n_0_0_38), .B2(res[10]), 
      .ZN(n_0_0_49));
   INV_X1 i_0_0_74 (.A(n_0_0_49), .ZN(n_0_245));
   AOI22_X1 i_0_0_75 (.A1(n_0_105), .A2(n_0_182), .B1(n_0_0_38), .B2(res[11]), 
      .ZN(n_0_0_50));
   INV_X1 i_0_0_76 (.A(n_0_0_50), .ZN(n_0_246));
   AOI22_X1 i_0_0_77 (.A1(n_0_105), .A2(n_0_183), .B1(n_0_0_38), .B2(res[12]), 
      .ZN(n_0_0_51));
   INV_X1 i_0_0_78 (.A(n_0_0_51), .ZN(n_0_247));
   AOI22_X1 i_0_0_79 (.A1(n_0_105), .A2(n_0_184), .B1(n_0_0_38), .B2(res[13]), 
      .ZN(n_0_0_52));
   INV_X1 i_0_0_80 (.A(n_0_0_52), .ZN(n_0_248));
   AOI22_X1 i_0_0_81 (.A1(n_0_105), .A2(n_0_185), .B1(n_0_0_38), .B2(res[14]), 
      .ZN(n_0_0_53));
   INV_X1 i_0_0_82 (.A(n_0_0_53), .ZN(n_0_249));
   AOI22_X1 i_0_0_83 (.A1(n_0_105), .A2(n_0_186), .B1(n_0_0_38), .B2(res[15]), 
      .ZN(n_0_0_54));
   INV_X1 i_0_0_84 (.A(n_0_0_54), .ZN(n_0_250));
   AOI22_X1 i_0_0_85 (.A1(n_0_105), .A2(n_0_187), .B1(n_0_0_38), .B2(res[16]), 
      .ZN(n_0_0_55));
   INV_X1 i_0_0_86 (.A(n_0_0_55), .ZN(n_0_251));
   AOI22_X1 i_0_0_87 (.A1(n_0_105), .A2(n_0_188), .B1(n_0_0_38), .B2(res[17]), 
      .ZN(n_0_0_56));
   INV_X1 i_0_0_88 (.A(n_0_0_56), .ZN(n_0_252));
   AOI22_X1 i_0_0_89 (.A1(n_0_105), .A2(n_0_189), .B1(n_0_0_38), .B2(res[18]), 
      .ZN(n_0_0_57));
   INV_X1 i_0_0_90 (.A(n_0_0_57), .ZN(n_0_253));
   AOI22_X1 i_0_0_91 (.A1(n_0_105), .A2(n_0_190), .B1(n_0_0_38), .B2(res[19]), 
      .ZN(n_0_0_58));
   INV_X1 i_0_0_92 (.A(n_0_0_58), .ZN(n_0_254));
   AOI22_X1 i_0_0_93 (.A1(n_0_105), .A2(n_0_191), .B1(n_0_0_38), .B2(res[20]), 
      .ZN(n_0_0_59));
   INV_X1 i_0_0_94 (.A(n_0_0_59), .ZN(n_0_255));
   AOI22_X1 i_0_0_95 (.A1(n_0_105), .A2(n_0_192), .B1(n_0_0_38), .B2(res[21]), 
      .ZN(n_0_0_60));
   INV_X1 i_0_0_96 (.A(n_0_0_60), .ZN(n_0_256));
   AOI22_X1 i_0_0_97 (.A1(n_0_105), .A2(n_0_193), .B1(n_0_0_38), .B2(res[22]), 
      .ZN(n_0_0_61));
   INV_X1 i_0_0_98 (.A(n_0_0_61), .ZN(n_0_257));
   AOI22_X1 i_0_0_99 (.A1(n_0_105), .A2(n_0_194), .B1(n_0_0_38), .B2(res[23]), 
      .ZN(n_0_0_62));
   INV_X1 i_0_0_100 (.A(n_0_0_62), .ZN(n_0_258));
   AOI22_X1 i_0_0_101 (.A1(n_0_105), .A2(n_0_195), .B1(n_0_0_38), .B2(res[24]), 
      .ZN(n_0_0_63));
   INV_X1 i_0_0_102 (.A(n_0_0_63), .ZN(n_0_259));
   AOI22_X1 i_0_0_103 (.A1(n_0_105), .A2(n_0_196), .B1(n_0_0_38), .B2(res[25]), 
      .ZN(n_0_0_64));
   INV_X1 i_0_0_104 (.A(n_0_0_64), .ZN(n_0_260));
   AOI22_X1 i_0_0_105 (.A1(n_0_105), .A2(n_0_197), .B1(n_0_0_38), .B2(res[26]), 
      .ZN(n_0_0_65));
   INV_X1 i_0_0_106 (.A(n_0_0_65), .ZN(n_0_261));
   AOI22_X1 i_0_0_107 (.A1(n_0_105), .A2(n_0_198), .B1(n_0_0_38), .B2(res[27]), 
      .ZN(n_0_0_66));
   INV_X1 i_0_0_108 (.A(n_0_0_66), .ZN(n_0_262));
   AOI22_X1 i_0_0_109 (.A1(n_0_105), .A2(n_0_199), .B1(n_0_0_38), .B2(res[28]), 
      .ZN(n_0_0_67));
   INV_X1 i_0_0_110 (.A(n_0_0_67), .ZN(n_0_263));
   AOI22_X1 i_0_0_111 (.A1(n_0_105), .A2(n_0_200), .B1(n_0_0_38), .B2(res[29]), 
      .ZN(n_0_0_68));
   INV_X1 i_0_0_112 (.A(n_0_0_68), .ZN(n_0_264));
   AOI22_X1 i_0_0_113 (.A1(n_0_105), .A2(n_0_201), .B1(n_0_0_38), .B2(res[30]), 
      .ZN(n_0_0_69));
   INV_X1 i_0_0_114 (.A(n_0_0_69), .ZN(n_0_265));
   AOI22_X1 i_0_0_115 (.A1(n_0_105), .A2(n_0_202), .B1(n_0_0_38), .B2(res[31]), 
      .ZN(n_0_0_70));
   INV_X1 i_0_0_116 (.A(n_0_0_70), .ZN(n_0_266));
   AOI22_X1 i_0_0_117 (.A1(n_0_105), .A2(n_0_203), .B1(n_0_0_38), .B2(res[32]), 
      .ZN(n_0_0_71));
   INV_X1 i_0_0_118 (.A(n_0_0_71), .ZN(n_0_267));
   AOI22_X1 i_0_0_119 (.A1(n_0_105), .A2(n_0_204), .B1(n_0_0_38), .B2(res[33]), 
      .ZN(n_0_0_72));
   INV_X1 i_0_0_120 (.A(n_0_0_72), .ZN(n_0_268));
   AOI22_X1 i_0_0_121 (.A1(n_0_105), .A2(n_0_205), .B1(n_0_0_38), .B2(res[34]), 
      .ZN(n_0_0_73));
   INV_X1 i_0_0_122 (.A(n_0_0_73), .ZN(n_0_269));
   AOI22_X1 i_0_0_123 (.A1(n_0_105), .A2(n_0_206), .B1(n_0_0_38), .B2(res[35]), 
      .ZN(n_0_0_74));
   INV_X1 i_0_0_124 (.A(n_0_0_74), .ZN(n_0_76));
   AOI22_X1 i_0_0_125 (.A1(n_0_105), .A2(n_0_207), .B1(n_0_0_38), .B2(res[36]), 
      .ZN(n_0_0_75));
   INV_X1 i_0_0_126 (.A(n_0_0_75), .ZN(n_0_77));
   AOI22_X1 i_0_0_127 (.A1(n_0_105), .A2(n_0_208), .B1(n_0_0_38), .B2(res[37]), 
      .ZN(n_0_0_76));
   INV_X1 i_0_0_128 (.A(n_0_0_76), .ZN(n_0_78));
   AOI22_X1 i_0_0_129 (.A1(n_0_105), .A2(n_0_209), .B1(n_0_0_38), .B2(res[38]), 
      .ZN(n_0_0_77));
   INV_X1 i_0_0_130 (.A(n_0_0_77), .ZN(n_0_79));
   AOI22_X1 i_0_0_131 (.A1(n_0_105), .A2(n_0_210), .B1(n_0_0_38), .B2(res[39]), 
      .ZN(n_0_0_78));
   INV_X1 i_0_0_132 (.A(n_0_0_78), .ZN(n_0_80));
   AOI22_X1 i_0_0_133 (.A1(n_0_105), .A2(n_0_211), .B1(n_0_0_38), .B2(res[40]), 
      .ZN(n_0_0_79));
   INV_X1 i_0_0_134 (.A(n_0_0_79), .ZN(n_0_81));
   AOI22_X1 i_0_0_135 (.A1(n_0_105), .A2(n_0_212), .B1(n_0_0_38), .B2(res[41]), 
      .ZN(n_0_0_80));
   INV_X1 i_0_0_136 (.A(n_0_0_80), .ZN(n_0_82));
   AOI22_X1 i_0_0_137 (.A1(n_0_105), .A2(n_0_213), .B1(n_0_0_38), .B2(res[42]), 
      .ZN(n_0_0_81));
   INV_X1 i_0_0_138 (.A(n_0_0_81), .ZN(n_0_83));
   AOI22_X1 i_0_0_139 (.A1(n_0_105), .A2(n_0_214), .B1(n_0_0_38), .B2(res[43]), 
      .ZN(n_0_0_82));
   INV_X1 i_0_0_140 (.A(n_0_0_82), .ZN(n_0_84));
   AOI22_X1 i_0_0_141 (.A1(n_0_105), .A2(n_0_215), .B1(n_0_0_38), .B2(res[44]), 
      .ZN(n_0_0_83));
   INV_X1 i_0_0_142 (.A(n_0_0_83), .ZN(n_0_85));
   AOI22_X1 i_0_0_143 (.A1(n_0_105), .A2(n_0_216), .B1(n_0_0_38), .B2(res[45]), 
      .ZN(n_0_0_84));
   INV_X1 i_0_0_144 (.A(n_0_0_84), .ZN(n_0_86));
   AOI22_X1 i_0_0_145 (.A1(n_0_105), .A2(n_0_217), .B1(n_0_0_38), .B2(res[46]), 
      .ZN(n_0_0_85));
   INV_X1 i_0_0_146 (.A(n_0_0_85), .ZN(n_0_87));
   AOI22_X1 i_0_0_147 (.A1(n_0_105), .A2(n_0_218), .B1(n_0_0_38), .B2(res[47]), 
      .ZN(n_0_0_86));
   INV_X1 i_0_0_148 (.A(n_0_0_86), .ZN(n_0_88));
   AOI22_X1 i_0_0_149 (.A1(n_0_105), .A2(n_0_219), .B1(n_0_0_38), .B2(res[48]), 
      .ZN(n_0_0_87));
   INV_X1 i_0_0_150 (.A(n_0_0_87), .ZN(n_0_89));
   AOI22_X1 i_0_0_151 (.A1(n_0_105), .A2(n_0_220), .B1(n_0_0_38), .B2(res[49]), 
      .ZN(n_0_0_88));
   INV_X1 i_0_0_152 (.A(n_0_0_88), .ZN(n_0_90));
   AOI22_X1 i_0_0_153 (.A1(n_0_105), .A2(n_0_221), .B1(n_0_0_38), .B2(res[50]), 
      .ZN(n_0_0_89));
   INV_X1 i_0_0_154 (.A(n_0_0_89), .ZN(n_0_91));
   AOI22_X1 i_0_0_155 (.A1(n_0_105), .A2(n_0_222), .B1(n_0_0_38), .B2(res[51]), 
      .ZN(n_0_0_90));
   INV_X1 i_0_0_156 (.A(n_0_0_90), .ZN(n_0_92));
   AOI22_X1 i_0_0_157 (.A1(n_0_105), .A2(n_0_223), .B1(n_0_0_38), .B2(res[52]), 
      .ZN(n_0_0_91));
   INV_X1 i_0_0_158 (.A(n_0_0_91), .ZN(n_0_93));
   AOI22_X1 i_0_0_159 (.A1(n_0_105), .A2(n_0_224), .B1(n_0_0_38), .B2(res[53]), 
      .ZN(n_0_0_92));
   INV_X1 i_0_0_160 (.A(n_0_0_92), .ZN(n_0_94));
   AOI22_X1 i_0_0_161 (.A1(n_0_105), .A2(n_0_225), .B1(n_0_0_38), .B2(res[54]), 
      .ZN(n_0_0_93));
   INV_X1 i_0_0_162 (.A(n_0_0_93), .ZN(n_0_95));
   AOI22_X1 i_0_0_163 (.A1(n_0_105), .A2(n_0_226), .B1(n_0_0_38), .B2(res[55]), 
      .ZN(n_0_0_94));
   INV_X1 i_0_0_164 (.A(n_0_0_94), .ZN(n_0_96));
   AOI22_X1 i_0_0_165 (.A1(n_0_105), .A2(n_0_227), .B1(n_0_0_38), .B2(res[56]), 
      .ZN(n_0_0_95));
   INV_X1 i_0_0_166 (.A(n_0_0_95), .ZN(n_0_97));
   AOI22_X1 i_0_0_167 (.A1(n_0_105), .A2(n_0_228), .B1(n_0_0_38), .B2(res[57]), 
      .ZN(n_0_0_96));
   INV_X1 i_0_0_168 (.A(n_0_0_96), .ZN(n_0_98));
   AOI22_X1 i_0_0_169 (.A1(n_0_105), .A2(n_0_229), .B1(n_0_0_38), .B2(res[58]), 
      .ZN(n_0_0_97));
   INV_X1 i_0_0_170 (.A(n_0_0_97), .ZN(n_0_99));
   AOI22_X1 i_0_0_171 (.A1(n_0_105), .A2(n_0_230), .B1(n_0_0_38), .B2(res[59]), 
      .ZN(n_0_0_98));
   INV_X1 i_0_0_172 (.A(n_0_0_98), .ZN(n_0_100));
   AOI22_X1 i_0_0_173 (.A1(n_0_105), .A2(n_0_231), .B1(n_0_0_38), .B2(res[60]), 
      .ZN(n_0_0_99));
   INV_X1 i_0_0_174 (.A(n_0_0_99), .ZN(n_0_101));
   AOI22_X1 i_0_0_175 (.A1(n_0_105), .A2(n_0_232), .B1(n_0_0_38), .B2(res[61]), 
      .ZN(n_0_0_100));
   INV_X1 i_0_0_176 (.A(n_0_0_100), .ZN(n_0_102));
   AOI22_X1 i_0_0_177 (.A1(n_0_105), .A2(n_0_233), .B1(n_0_0_38), .B2(res[62]), 
      .ZN(n_0_0_101));
   INV_X1 i_0_0_178 (.A(n_0_0_101), .ZN(n_0_103));
   AOI22_X1 i_0_0_179 (.A1(n_0_105), .A2(n_0_234), .B1(n_0_0_38), .B2(res[63]), 
      .ZN(n_0_0_102));
   INV_X1 i_0_0_180 (.A(n_0_0_102), .ZN(n_0_104));
   INV_X1 i_0_0_181 (.A(i[4]), .ZN(n_0_0_103));
   AND2_X1 i_0_0_182 (.A1(n_0_0_103), .A2(i[3]), .ZN(n_0_0_104));
   NOR2_X1 i_0_0_183 (.A1(n_0_0_103), .A2(i[3]), .ZN(n_0_0_105));
   AOI22_X1 i_0_0_184 (.A1(n_0_0_104), .A2(read_data[11]), .B1(n_0_0_105), 
      .B2(read_data[19]), .ZN(n_0_0_106));
   NAND2_X1 i_0_0_185 (.A1(i[4]), .A2(i[3]), .ZN(n_0_0_107));
   INV_X1 i_0_0_186 (.A(n_0_0_107), .ZN(n_0_0_108));
   AOI22_X1 i_0_0_187 (.A1(n_0_0_108), .A2(read_data[27]), .B1(n_0_0_35), 
      .B2(read_data[3]), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_106), .A2(n_0_0_109), .ZN(n_0_0_110));
   INV_X1 i_0_0_189 (.A(n_0_0_110), .ZN(n_0_0_111));
   AOI22_X1 i_0_0_190 (.A1(n_0_0_104), .A2(read_data[14]), .B1(n_0_0_105), 
      .B2(read_data[22]), .ZN(n_0_0_112));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_108), .A2(read_data[30]), .B1(n_0_0_35), 
      .B2(read_data[6]), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_192 (.A1(n_0_0_112), .A2(n_0_0_113), .ZN(n_0_0_114));
   INV_X1 i_0_0_193 (.A(n_0_0_114), .ZN(n_0_0_115));
   OAI33_X1 i_0_0_194 (.A1(n_0_0_111), .A2(i[1]), .A3(i[0]), .B1(n_0_0_115), 
      .B2(n_0_0_6), .B3(n_0_0_1), .ZN(n_0_0_116));
   NAND3_X1 i_0_0_195 (.A1(n_0_0_116), .A2(n_0_0_17), .A3(i[2]), .ZN(n_0_0_117));
   INV_X1 i_0_0_196 (.A(read_data[31]), .ZN(n_0_0_118));
   NOR3_X1 i_0_0_197 (.A1(n_0_0_36), .A2(n_0_0_17), .A3(n_0_0_118), .ZN(
      n_0_0_119));
   AOI222_X1 i_0_0_198 (.A1(n_0_0_108), .A2(read_data[24]), .B1(n_0_0_104), 
      .B2(read_data[8]), .C1(n_0_0_105), .C2(read_data[16]), .ZN(n_0_0_120));
   INV_X1 i_0_0_199 (.A(n_0_0_120), .ZN(n_0_0_121));
   AOI21_X1 i_0_0_200 (.A(n_0_0_121), .B1(read_data[0]), .B2(n_0_0_35), .ZN(
      n_0_0_122));
   NOR2_X1 i_0_0_201 (.A1(i[5]), .A2(i[1]), .ZN(n_0_0_123));
   NAND3_X1 i_0_0_202 (.A1(n_0_0_123), .A2(i[0]), .A3(n_0_0_7), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_203 (.A1(n_0_0_104), .A2(read_data[9]), .B1(n_0_0_105), 
      .B2(read_data[17]), .ZN(n_0_0_125));
   AOI22_X1 i_0_0_204 (.A1(n_0_0_108), .A2(read_data[25]), .B1(n_0_0_35), 
      .B2(read_data[1]), .ZN(n_0_0_126));
   NAND2_X1 i_0_0_205 (.A1(n_0_0_125), .A2(n_0_0_126), .ZN(n_0_0_127));
   INV_X1 i_0_0_206 (.A(n_0_0_127), .ZN(n_0_0_128));
   INV_X1 i_0_0_207 (.A(n_0_0_34), .ZN(n_0_0_129));
   NAND2_X1 i_0_0_208 (.A1(n_0_0_17), .A2(i[1]), .ZN(n_0_0_130));
   OR2_X1 i_0_0_209 (.A1(n_0_0_129), .A2(n_0_0_130), .ZN(n_0_0_131));
   OAI22_X1 i_0_0_210 (.A1(n_0_0_122), .A2(n_0_0_124), .B1(n_0_0_128), .B2(
      n_0_0_131), .ZN(n_0_0_132));
   AOI222_X1 i_0_0_211 (.A1(n_0_0_108), .A2(read_data[23]), .B1(n_0_0_105), 
      .B2(read_data[15]), .C1(n_0_0_104), .C2(read_data[7]), .ZN(n_0_0_133));
   AOI22_X1 i_0_0_212 (.A1(n_0_0_104), .A2(read_data[12]), .B1(n_0_0_105), 
      .B2(read_data[20]), .ZN(n_0_0_134));
   AOI22_X1 i_0_0_213 (.A1(n_0_0_108), .A2(read_data[28]), .B1(n_0_0_35), 
      .B2(read_data[4]), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_214 (.A1(n_0_0_134), .A2(n_0_0_135), .ZN(n_0_0_136));
   INV_X1 i_0_0_215 (.A(n_0_0_136), .ZN(n_0_0_137));
   NAND2_X1 i_0_0_216 (.A1(i[0]), .A2(i[2]), .ZN(n_0_0_138));
   OAI22_X1 i_0_0_217 (.A1(n_0_0_133), .A2(n_0_0_129), .B1(n_0_0_137), .B2(
      n_0_0_138), .ZN(n_0_0_139));
   AOI211_X1 i_0_0_218 (.A(n_0_0_119), .B(n_0_0_132), .C1(n_0_0_123), .C2(
      n_0_0_139), .ZN(n_0_0_140));
   AOI22_X1 i_0_0_219 (.A1(n_0_0_104), .A2(read_data[13]), .B1(n_0_0_105), 
      .B2(read_data[21]), .ZN(n_0_0_141));
   AOI22_X1 i_0_0_220 (.A1(n_0_0_108), .A2(read_data[29]), .B1(n_0_0_35), 
      .B2(read_data[5]), .ZN(n_0_0_142));
   NAND2_X1 i_0_0_221 (.A1(n_0_0_141), .A2(n_0_0_142), .ZN(n_0_0_143));
   NOR2_X1 i_0_0_222 (.A1(n_0_0_7), .A2(i[0]), .ZN(n_0_0_144));
   AOI22_X1 i_0_0_223 (.A1(n_0_0_104), .A2(read_data[10]), .B1(n_0_0_105), 
      .B2(read_data[18]), .ZN(n_0_0_145));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_108), .A2(read_data[26]), .B1(n_0_0_35), 
      .B2(read_data[2]), .ZN(n_0_0_146));
   NAND2_X1 i_0_0_225 (.A1(n_0_0_145), .A2(n_0_0_146), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_226 (.A1(n_0_0_7), .A2(i[0]), .ZN(n_0_0_148));
   INV_X1 i_0_0_227 (.A(n_0_0_148), .ZN(n_0_0_149));
   AOI22_X1 i_0_0_228 (.A1(n_0_0_143), .A2(n_0_0_144), .B1(n_0_0_147), .B2(
      n_0_0_149), .ZN(n_0_0_150));
   OAI211_X1 i_0_0_229 (.A(n_0_0_117), .B(n_0_0_140), .C1(n_0_0_130), .C2(
      n_0_0_150), .ZN(n_0_0_151));
   INV_X1 i_0_0_230 (.A(n_0_0_147), .ZN(n_0_0_152));
   INV_X1 i_0_0_231 (.A(n_0_0_143), .ZN(n_0_0_153));
   OAI33_X1 i_0_0_232 (.A1(n_0_0_152), .A2(i[1]), .A3(i[0]), .B1(n_0_0_153), 
      .B2(n_0_0_6), .B3(n_0_0_1), .ZN(n_0_0_154));
   NAND3_X1 i_0_0_233 (.A1(n_0_0_154), .A2(n_0_0_17), .A3(i[2]), .ZN(n_0_0_155));
   AOI222_X1 i_0_0_234 (.A1(read_data[22]), .A2(n_0_0_108), .B1(n_0_0_105), 
      .B2(read_data[14]), .C1(n_0_0_104), .C2(read_data[6]), .ZN(n_0_0_156));
   OAI22_X1 i_0_0_235 (.A1(n_0_0_156), .A2(n_0_0_129), .B1(n_0_0_111), .B2(
      n_0_0_138), .ZN(n_0_0_157));
   INV_X1 i_0_0_236 (.A(read_data[30]), .ZN(n_0_0_158));
   OAI22_X1 i_0_0_237 (.A1(n_0_0_129), .A2(n_0_0_158), .B1(n_0_0_148), .B2(
      n_0_0_118), .ZN(n_0_0_159));
   INV_X1 i_0_0_238 (.A(n_0_0_35), .ZN(n_0_0_160));
   NOR3_X1 i_0_0_239 (.A1(n_0_0_160), .A2(n_0_0_17), .A3(i[1]), .ZN(n_0_0_161));
   AOI22_X1 i_0_0_240 (.A1(n_0_0_157), .A2(n_0_0_123), .B1(n_0_0_159), .B2(
      n_0_0_161), .ZN(n_0_0_162));
   AOI22_X1 i_0_0_241 (.A1(n_0_0_127), .A2(n_0_0_149), .B1(n_0_0_136), .B2(
      n_0_0_144), .ZN(n_0_0_163));
   OAI211_X1 i_0_0_242 (.A(n_0_0_155), .B(n_0_0_162), .C1(n_0_0_130), .C2(
      n_0_0_163), .ZN(n_0_0_164));
   OAI22_X1 i_0_0_243 (.A1(n_0_0_122), .A2(n_0_0_131), .B1(n_0_0_124), .B2(
      n_0_0_133), .ZN(n_0_0_165));
   NOR2_X1 i_0_0_244 (.A1(n_0_0_164), .A2(n_0_0_165), .ZN(n_0_0_166));
   INV_X1 i_0_0_245 (.A(n_0_0_166), .ZN(n_0_0_167));
   INV_X1 i_0_0_246 (.A(n_0_0_151), .ZN(n_0_0_168));
   OAI22_X1 i_0_0_247 (.A1(n_0_0_151), .A2(n_0_0_167), .B1(n_0_0_168), .B2(
      n_0_0_166), .ZN(n_0_0_169));
   INV_X1 i_0_0_248 (.A(read_data2[0]), .ZN(n_0_0_170));
   OR2_X1 i_0_0_249 (.A1(n_0_0_169), .A2(n_0_0_170), .ZN(n_0_0_171));
   NOR2_X1 i_0_0_250 (.A1(shift[5]), .A2(shift[3]), .ZN(n_0_0_172));
   INV_X1 i_0_0_251 (.A(shift[4]), .ZN(n_0_0_173));
   NAND3_X1 i_0_0_252 (.A1(n_0_0_172), .A2(n_0_0_173), .A3(n_0_0_23), .ZN(
      n_0_0_174));
   NOR2_X1 i_0_0_253 (.A1(n_0_0_174), .A2(shift[1]), .ZN(n_0_0_175));
   INV_X1 i_0_0_254 (.A(n_0_0_175), .ZN(n_0_0_176));
   NOR3_X1 i_0_0_255 (.A1(n_0_0_171), .A2(shift[0]), .A3(n_0_0_176), .ZN(n_0_108));
   INV_X1 i_0_0_256 (.A(read_data[0]), .ZN(n_0_0_177));
   NOR3_X1 i_0_0_257 (.A1(n_0_0_36), .A2(i[5]), .A3(n_0_0_177), .ZN(n_0_0_178));
   INV_X1 i_0_0_258 (.A(n_0_0_124), .ZN(n_0_0_179));
   INV_X1 i_0_0_259 (.A(n_0_0_131), .ZN(n_0_0_180));
   AOI221_X1 i_0_0_260 (.A(n_0_0_178), .B1(n_0_0_127), .B2(n_0_0_179), .C1(
      n_0_0_180), .C2(n_0_0_147), .ZN(n_0_0_181));
   AOI22_X1 i_0_0_261 (.A1(n_0_0_110), .A2(n_0_0_149), .B1(n_0_0_114), .B2(
      n_0_0_144), .ZN(n_0_0_182));
   OAI21_X1 i_0_0_262 (.A(n_0_0_181), .B1(n_0_0_130), .B2(n_0_0_182), .ZN(
      n_0_0_183));
   INV_X1 i_0_0_263 (.A(read_data[7]), .ZN(n_0_0_184));
   OAI22_X1 i_0_0_264 (.A1(n_0_0_160), .A2(n_0_0_184), .B1(n_0_0_107), .B2(
      n_0_0_118), .ZN(n_0_0_185));
   AOI221_X1 i_0_0_265 (.A(n_0_0_185), .B1(read_data[23]), .B2(n_0_0_105), 
      .C1(read_data[15]), .C2(n_0_0_104), .ZN(n_0_0_186));
   OAI33_X1 i_0_0_266 (.A1(n_0_0_186), .A2(n_0_0_6), .A3(n_0_0_1), .B1(n_0_0_137), 
      .B2(i[1]), .B3(i[0]), .ZN(n_0_0_187));
   AND3_X1 i_0_0_267 (.A1(n_0_0_187), .A2(n_0_0_17), .A3(i[2]), .ZN(n_0_0_188));
   OAI22_X1 i_0_0_268 (.A1(n_0_0_120), .A2(n_0_0_129), .B1(n_0_0_153), .B2(
      n_0_0_138), .ZN(n_0_0_189));
   AOI211_X1 i_0_0_269 (.A(n_0_0_183), .B(n_0_0_188), .C1(n_0_0_123), .C2(
      n_0_0_189), .ZN(n_0_0_190));
   INV_X1 i_0_0_270 (.A(n_0_0_190), .ZN(n_0_0_191));
   NOR3_X1 i_0_0_271 (.A1(n_0_0_168), .A2(n_0_0_166), .A3(n_0_0_191), .ZN(
      n_0_0_192));
   INV_X1 i_0_0_272 (.A(n_0_0_192), .ZN(n_0_0_193));
   NAND3_X1 i_0_0_273 (.A1(n_0_0_168), .A2(n_0_0_166), .A3(n_0_0_191), .ZN(
      n_0_0_194));
   AOI21_X1 i_0_0_274 (.A(n_0_0_170), .B1(n_0_0_193), .B2(n_0_0_194), .ZN(
      n_0_0_195));
   NOR2_X1 i_0_0_275 (.A1(n_0_0_169), .A2(n_0_0_190), .ZN(n_0_0_196));
   NOR2_X1 i_0_0_276 (.A1(n_0_0_169), .A2(n_0_0_191), .ZN(n_0_0_197));
   AOI221_X1 i_0_0_277 (.A(n_0_0_195), .B1(n_0_0_196), .B2(n_0_4), .C1(
      read_data2[1]), .C2(n_0_0_197), .ZN(n_0_0_198));
   OAI33_X1 i_0_0_278 (.A1(n_0_0_198), .A2(shift[0]), .A3(n_0_0_176), .B1(
      n_0_0_171), .B2(n_0_0_19), .B3(n_0_0_176), .ZN(n_0_109));
   NAND2_X1 i_0_0_279 (.A1(n_0_0_175), .A2(shift[0]), .ZN(n_0_0_199));
   INV_X1 i_0_0_280 (.A(n_0_0_194), .ZN(n_0_0_200));
   AOI22_X1 i_0_0_281 (.A1(n_0_0_197), .A2(read_data2[2]), .B1(n_0_0_200), 
      .B2(n_0_35), .ZN(n_0_0_201));
   AOI22_X1 i_0_0_282 (.A1(n_0_0_196), .A2(n_0_5), .B1(read_data2[1]), .B2(
      n_0_0_192), .ZN(n_0_0_202));
   NAND2_X1 i_0_0_283 (.A1(n_0_0_201), .A2(n_0_0_202), .ZN(n_0_0_203));
   INV_X1 i_0_0_284 (.A(n_0_0_171), .ZN(n_0_0_204));
   NOR2_X1 i_0_0_285 (.A1(n_0_0_174), .A2(n_0_0_24), .ZN(n_0_0_205));
   AOI22_X1 i_0_0_286 (.A1(n_0_0_203), .A2(n_0_0_175), .B1(n_0_0_204), .B2(
      n_0_0_205), .ZN(n_0_0_206));
   OAI22_X1 i_0_0_287 (.A1(n_0_0_198), .A2(n_0_0_199), .B1(n_0_0_206), .B2(
      shift[0]), .ZN(n_0_110));
   AOI22_X1 i_0_0_288 (.A1(n_0_0_197), .A2(read_data2[3]), .B1(n_0_0_200), 
      .B2(n_0_36), .ZN(n_0_0_207));
   AOI22_X1 i_0_0_289 (.A1(n_0_0_196), .A2(n_0_6), .B1(read_data2[2]), .B2(
      n_0_0_192), .ZN(n_0_0_208));
   NAND2_X1 i_0_0_290 (.A1(n_0_0_207), .A2(n_0_0_208), .ZN(n_0_0_209));
   INV_X1 i_0_0_291 (.A(n_0_0_198), .ZN(n_0_0_210));
   AOI22_X1 i_0_0_292 (.A1(n_0_0_175), .A2(n_0_0_209), .B1(n_0_0_210), .B2(
      n_0_0_205), .ZN(n_0_0_211));
   AOI22_X1 i_0_0_293 (.A1(n_0_0_211), .A2(n_0_0_19), .B1(n_0_0_206), .B2(
      shift[0]), .ZN(n_0_111));
   AOI22_X1 i_0_0_294 (.A1(n_0_0_197), .A2(read_data2[4]), .B1(n_0_0_200), 
      .B2(n_0_37), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_295 (.A1(n_0_0_196), .A2(n_0_7), .B1(read_data2[3]), .B2(
      n_0_0_192), .ZN(n_0_0_213));
   NAND2_X1 i_0_0_296 (.A1(n_0_0_212), .A2(n_0_0_213), .ZN(n_0_0_214));
   INV_X1 i_0_0_297 (.A(n_0_0_214), .ZN(n_0_0_215));
   NAND3_X1 i_0_0_298 (.A1(n_0_0_172), .A2(n_0_0_173), .A3(shift[2]), .ZN(
      n_0_0_216));
   OAI22_X1 i_0_0_299 (.A1(n_0_0_215), .A2(n_0_0_174), .B1(n_0_0_171), .B2(
      n_0_0_216), .ZN(n_0_0_217));
   AOI22_X1 i_0_0_300 (.A1(n_0_0_217), .A2(n_0_0_24), .B1(n_0_0_203), .B2(
      n_0_0_205), .ZN(n_0_0_218));
   OAI22_X1 i_0_0_301 (.A1(n_0_0_218), .A2(shift[0]), .B1(n_0_0_19), .B2(
      n_0_0_211), .ZN(n_0_112));
   AOI22_X1 i_0_0_302 (.A1(n_0_0_197), .A2(read_data2[5]), .B1(n_0_0_200), 
      .B2(n_0_38), .ZN(n_0_0_219));
   AOI22_X1 i_0_0_303 (.A1(n_0_0_196), .A2(n_0_8), .B1(read_data2[4]), .B2(
      n_0_0_192), .ZN(n_0_0_220));
   NAND2_X1 i_0_0_304 (.A1(n_0_0_219), .A2(n_0_0_220), .ZN(n_0_0_221));
   INV_X1 i_0_0_305 (.A(n_0_0_221), .ZN(n_0_0_222));
   OAI22_X1 i_0_0_306 (.A1(n_0_0_198), .A2(n_0_0_216), .B1(n_0_0_222), .B2(
      n_0_0_174), .ZN(n_0_0_223));
   AOI22_X1 i_0_0_307 (.A1(n_0_0_223), .A2(n_0_0_24), .B1(n_0_0_209), .B2(
      n_0_0_205), .ZN(n_0_0_224));
   OAI22_X1 i_0_0_308 (.A1(n_0_0_224), .A2(shift[0]), .B1(n_0_0_218), .B2(
      n_0_0_19), .ZN(n_0_113));
   INV_X1 i_0_0_309 (.A(n_0_0_203), .ZN(n_0_0_225));
   AOI22_X1 i_0_0_310 (.A1(n_0_0_196), .A2(n_0_9), .B1(n_0_0_200), .B2(n_0_39), 
      .ZN(n_0_0_226));
   AOI22_X1 i_0_0_311 (.A1(n_0_0_197), .A2(read_data2[6]), .B1(read_data2[5]), 
      .B2(n_0_0_192), .ZN(n_0_0_227));
   NAND2_X1 i_0_0_312 (.A1(n_0_0_226), .A2(n_0_0_227), .ZN(n_0_0_228));
   INV_X1 i_0_0_313 (.A(n_0_0_228), .ZN(n_0_0_229));
   OAI22_X1 i_0_0_314 (.A1(n_0_0_225), .A2(n_0_0_216), .B1(n_0_0_229), .B2(
      n_0_0_174), .ZN(n_0_0_230));
   OAI22_X1 i_0_0_315 (.A1(n_0_0_230), .A2(shift[1]), .B1(n_0_0_217), .B2(
      n_0_0_24), .ZN(n_0_0_231));
   OAI22_X1 i_0_0_316 (.A1(n_0_0_224), .A2(n_0_0_19), .B1(n_0_0_231), .B2(
      shift[0]), .ZN(n_0_114));
   AOI22_X1 i_0_0_317 (.A1(n_0_0_197), .A2(read_data2[7]), .B1(n_0_0_200), 
      .B2(n_0_40), .ZN(n_0_0_232));
   AOI22_X1 i_0_0_318 (.A1(n_0_0_196), .A2(n_0_10), .B1(read_data2[6]), .B2(
      n_0_0_192), .ZN(n_0_0_233));
   NAND2_X1 i_0_0_319 (.A1(n_0_0_232), .A2(n_0_0_233), .ZN(n_0_0_234));
   INV_X1 i_0_0_320 (.A(n_0_0_234), .ZN(n_0_0_235));
   INV_X1 i_0_0_321 (.A(n_0_0_209), .ZN(n_0_0_236));
   OAI22_X1 i_0_0_322 (.A1(n_0_0_235), .A2(n_0_0_174), .B1(n_0_0_236), .B2(
      n_0_0_216), .ZN(n_0_0_237));
   OAI22_X1 i_0_0_323 (.A1(n_0_0_223), .A2(n_0_0_24), .B1(n_0_0_237), .B2(
      shift[1]), .ZN(n_0_0_238));
   OAI22_X1 i_0_0_324 (.A1(n_0_0_238), .A2(shift[0]), .B1(n_0_0_231), .B2(
      n_0_0_19), .ZN(n_0_115));
   AOI22_X1 i_0_0_325 (.A1(n_0_0_197), .A2(read_data2[8]), .B1(n_0_0_200), 
      .B2(n_0_41), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_326 (.A1(n_0_0_196), .A2(n_0_11), .B1(read_data2[7]), .B2(
      n_0_0_192), .ZN(n_0_0_240));
   NAND2_X1 i_0_0_327 (.A1(n_0_0_239), .A2(n_0_0_240), .ZN(n_0_0_241));
   AND2_X1 i_0_0_328 (.A1(n_0_0_172), .A2(n_0_0_173), .ZN(n_0_0_242));
   NAND2_X1 i_0_0_329 (.A1(n_0_0_33), .A2(shift[3]), .ZN(n_0_0_243));
   NOR2_X1 i_0_0_330 (.A1(n_0_0_243), .A2(shift[4]), .ZN(n_0_0_244));
   AOI22_X1 i_0_0_331 (.A1(n_0_0_241), .A2(n_0_0_242), .B1(n_0_0_204), .B2(
      n_0_0_244), .ZN(n_0_0_245));
   OAI22_X1 i_0_0_332 (.A1(n_0_0_245), .A2(shift[2]), .B1(n_0_0_215), .B2(
      n_0_0_216), .ZN(n_0_0_246));
   AOI22_X1 i_0_0_333 (.A1(n_0_0_246), .A2(n_0_0_24), .B1(n_0_0_230), .B2(
      shift[1]), .ZN(n_0_0_247));
   OAI22_X1 i_0_0_334 (.A1(n_0_0_238), .A2(n_0_0_19), .B1(n_0_0_247), .B2(
      shift[0]), .ZN(n_0_116));
   AOI22_X1 i_0_0_335 (.A1(n_0_0_197), .A2(read_data2[9]), .B1(n_0_0_200), 
      .B2(n_0_42), .ZN(n_0_0_248));
   AOI22_X1 i_0_0_336 (.A1(n_0_0_196), .A2(n_0_12), .B1(read_data2[8]), .B2(
      n_0_0_192), .ZN(n_0_0_249));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_248), .A2(n_0_0_249), .ZN(n_0_0_250));
   AOI22_X1 i_0_0_338 (.A1(n_0_0_242), .A2(n_0_0_250), .B1(n_0_0_210), .B2(
      n_0_0_244), .ZN(n_0_0_251));
   OAI22_X1 i_0_0_339 (.A1(n_0_0_251), .A2(shift[2]), .B1(n_0_0_222), .B2(
      n_0_0_216), .ZN(n_0_0_252));
   AOI22_X1 i_0_0_340 (.A1(n_0_0_252), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_237), .ZN(n_0_0_253));
   OAI22_X1 i_0_0_341 (.A1(n_0_0_253), .A2(shift[0]), .B1(n_0_0_247), .B2(
      n_0_0_19), .ZN(n_0_117));
   AOI22_X1 i_0_0_342 (.A1(n_0_0_196), .A2(n_0_13), .B1(n_0_0_200), .B2(n_0_43), 
      .ZN(n_0_0_254));
   AOI22_X1 i_0_0_343 (.A1(n_0_0_197), .A2(read_data2[10]), .B1(read_data2[9]), 
      .B2(n_0_0_192), .ZN(n_0_0_255));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_254), .A2(n_0_0_255), .ZN(n_0_0_256));
   AOI22_X1 i_0_0_345 (.A1(n_0_0_203), .A2(n_0_0_244), .B1(n_0_0_256), .B2(
      n_0_0_242), .ZN(n_0_0_257));
   OAI22_X1 i_0_0_346 (.A1(n_0_0_257), .A2(shift[2]), .B1(n_0_0_229), .B2(
      n_0_0_216), .ZN(n_0_0_258));
   AOI22_X1 i_0_0_347 (.A1(n_0_0_258), .A2(n_0_0_24), .B1(n_0_0_246), .B2(
      shift[1]), .ZN(n_0_0_259));
   OAI22_X1 i_0_0_348 (.A1(n_0_0_253), .A2(n_0_0_19), .B1(n_0_0_259), .B2(
      shift[0]), .ZN(n_0_118));
   AOI22_X1 i_0_0_349 (.A1(n_0_0_196), .A2(n_0_14), .B1(n_0_0_200), .B2(n_0_44), 
      .ZN(n_0_0_260));
   AOI22_X1 i_0_0_350 (.A1(n_0_0_197), .A2(read_data2[11]), .B1(read_data2[10]), 
      .B2(n_0_0_192), .ZN(n_0_0_261));
   NAND2_X1 i_0_0_351 (.A1(n_0_0_260), .A2(n_0_0_261), .ZN(n_0_0_262));
   AOI22_X1 i_0_0_352 (.A1(n_0_0_262), .A2(n_0_0_242), .B1(n_0_0_209), .B2(
      n_0_0_244), .ZN(n_0_0_263));
   OAI22_X1 i_0_0_353 (.A1(n_0_0_263), .A2(shift[2]), .B1(n_0_0_235), .B2(
      n_0_0_216), .ZN(n_0_0_264));
   AOI22_X1 i_0_0_354 (.A1(n_0_0_264), .A2(n_0_0_24), .B1(n_0_0_252), .B2(
      shift[1]), .ZN(n_0_0_265));
   OAI22_X1 i_0_0_355 (.A1(n_0_0_265), .A2(shift[0]), .B1(n_0_0_259), .B2(
      n_0_0_19), .ZN(n_0_119));
   AOI22_X1 i_0_0_356 (.A1(n_0_0_197), .A2(read_data2[12]), .B1(n_0_0_196), 
      .B2(n_0_15), .ZN(n_0_0_266));
   AOI22_X1 i_0_0_357 (.A1(n_0_0_200), .A2(n_0_45), .B1(read_data2[11]), 
      .B2(n_0_0_192), .ZN(n_0_0_267));
   NAND2_X1 i_0_0_358 (.A1(n_0_0_266), .A2(n_0_0_267), .ZN(n_0_0_268));
   AOI22_X1 i_0_0_359 (.A1(n_0_0_268), .A2(n_0_0_242), .B1(n_0_0_214), .B2(
      n_0_0_244), .ZN(n_0_0_269));
   OAI22_X1 i_0_0_360 (.A1(n_0_0_269), .A2(shift[2]), .B1(n_0_0_245), .B2(
      n_0_0_23), .ZN(n_0_0_270));
   AOI22_X1 i_0_0_361 (.A1(n_0_0_270), .A2(n_0_0_24), .B1(n_0_0_258), .B2(
      shift[1]), .ZN(n_0_0_271));
   OAI22_X1 i_0_0_362 (.A1(n_0_0_265), .A2(n_0_0_19), .B1(n_0_0_271), .B2(
      shift[0]), .ZN(n_0_120));
   AOI22_X1 i_0_0_363 (.A1(n_0_0_197), .A2(read_data2[13]), .B1(n_0_0_200), 
      .B2(n_0_46), .ZN(n_0_0_272));
   AOI22_X1 i_0_0_364 (.A1(n_0_0_196), .A2(n_0_16), .B1(read_data2[12]), 
      .B2(n_0_0_192), .ZN(n_0_0_273));
   NAND2_X1 i_0_0_365 (.A1(n_0_0_272), .A2(n_0_0_273), .ZN(n_0_0_274));
   AOI22_X1 i_0_0_366 (.A1(n_0_0_221), .A2(n_0_0_244), .B1(n_0_0_274), .B2(
      n_0_0_242), .ZN(n_0_0_275));
   OAI22_X1 i_0_0_367 (.A1(n_0_0_251), .A2(n_0_0_23), .B1(n_0_0_275), .B2(
      shift[2]), .ZN(n_0_0_276));
   AOI22_X1 i_0_0_368 (.A1(n_0_0_276), .A2(n_0_0_24), .B1(n_0_0_264), .B2(
      shift[1]), .ZN(n_0_0_277));
   OAI22_X1 i_0_0_369 (.A1(n_0_0_277), .A2(shift[0]), .B1(n_0_0_271), .B2(
      n_0_0_19), .ZN(n_0_121));
   AOI22_X1 i_0_0_370 (.A1(n_0_0_196), .A2(n_0_17), .B1(n_0_0_200), .B2(n_0_47), 
      .ZN(n_0_0_278));
   AOI22_X1 i_0_0_371 (.A1(n_0_0_197), .A2(read_data2[14]), .B1(read_data2[13]), 
      .B2(n_0_0_192), .ZN(n_0_0_279));
   NAND2_X1 i_0_0_372 (.A1(n_0_0_278), .A2(n_0_0_279), .ZN(n_0_0_280));
   AOI22_X1 i_0_0_373 (.A1(n_0_0_280), .A2(n_0_0_242), .B1(n_0_0_228), .B2(
      n_0_0_244), .ZN(n_0_0_281));
   OAI22_X1 i_0_0_374 (.A1(n_0_0_257), .A2(n_0_0_23), .B1(n_0_0_281), .B2(
      shift[2]), .ZN(n_0_0_282));
   AOI22_X1 i_0_0_375 (.A1(n_0_0_282), .A2(n_0_0_24), .B1(n_0_0_270), .B2(
      shift[1]), .ZN(n_0_0_283));
   OAI22_X1 i_0_0_376 (.A1(n_0_0_277), .A2(n_0_0_19), .B1(n_0_0_283), .B2(
      shift[0]), .ZN(n_0_122));
   AOI22_X1 i_0_0_377 (.A1(n_0_0_196), .A2(n_0_18), .B1(n_0_0_200), .B2(n_0_48), 
      .ZN(n_0_0_284));
   AOI22_X1 i_0_0_378 (.A1(n_0_0_197), .A2(read_data2[15]), .B1(read_data2[14]), 
      .B2(n_0_0_192), .ZN(n_0_0_285));
   NAND2_X1 i_0_0_379 (.A1(n_0_0_284), .A2(n_0_0_285), .ZN(n_0_0_286));
   AOI22_X1 i_0_0_380 (.A1(n_0_0_234), .A2(n_0_0_244), .B1(n_0_0_286), .B2(
      n_0_0_242), .ZN(n_0_0_287));
   AOI22_X1 i_0_0_381 (.A1(n_0_0_263), .A2(shift[2]), .B1(n_0_0_287), .B2(
      n_0_0_23), .ZN(n_0_0_288));
   AOI22_X1 i_0_0_382 (.A1(n_0_0_288), .A2(n_0_0_24), .B1(n_0_0_276), .B2(
      shift[1]), .ZN(n_0_0_289));
   OAI22_X1 i_0_0_383 (.A1(n_0_0_289), .A2(shift[0]), .B1(n_0_0_283), .B2(
      n_0_0_19), .ZN(n_0_123));
   AOI22_X1 i_0_0_384 (.A1(n_0_0_196), .A2(n_0_19), .B1(n_0_0_200), .B2(n_0_49), 
      .ZN(n_0_0_290));
   AOI22_X1 i_0_0_385 (.A1(n_0_0_197), .A2(read_data2[16]), .B1(read_data2[15]), 
      .B2(n_0_0_192), .ZN(n_0_0_291));
   NAND2_X1 i_0_0_386 (.A1(n_0_0_290), .A2(n_0_0_291), .ZN(n_0_0_292));
   AOI22_X1 i_0_0_387 (.A1(n_0_0_292), .A2(n_0_0_173), .B1(shift[4]), .B2(
      n_0_0_204), .ZN(n_0_0_293));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_293), .A2(shift[5]), .ZN(n_0_0_294));
   INV_X1 i_0_0_389 (.A(shift[3]), .ZN(n_0_0_295));
   AOI22_X1 i_0_0_390 (.A1(n_0_0_294), .A2(n_0_0_295), .B1(n_0_0_241), .B2(
      n_0_0_244), .ZN(n_0_0_296));
   OAI22_X1 i_0_0_391 (.A1(n_0_0_296), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_269), .ZN(n_0_0_297));
   AOI22_X1 i_0_0_392 (.A1(n_0_0_297), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_282), .ZN(n_0_0_298));
   OAI22_X1 i_0_0_393 (.A1(n_0_0_298), .A2(shift[0]), .B1(n_0_0_19), .B2(
      n_0_0_289), .ZN(n_0_124));
   AOI22_X1 i_0_0_394 (.A1(n_0_0_196), .A2(n_0_20), .B1(n_0_0_200), .B2(n_0_50), 
      .ZN(n_0_0_299));
   AOI22_X1 i_0_0_395 (.A1(n_0_0_197), .A2(read_data2[17]), .B1(read_data2[16]), 
      .B2(n_0_0_192), .ZN(n_0_0_300));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_299), .A2(n_0_0_300), .ZN(n_0_0_301));
   OAI22_X1 i_0_0_397 (.A1(n_0_0_301), .A2(shift[4]), .B1(n_0_0_210), .B2(
      n_0_0_173), .ZN(n_0_0_302));
   INV_X1 i_0_0_398 (.A(n_0_0_302), .ZN(n_0_0_303));
   AOI22_X1 i_0_0_399 (.A1(n_0_0_303), .A2(n_0_0_172), .B1(n_0_0_244), .B2(
      n_0_0_250), .ZN(n_0_0_304));
   OAI22_X1 i_0_0_400 (.A1(n_0_0_304), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_275), .ZN(n_0_0_305));
   AOI22_X1 i_0_0_401 (.A1(n_0_0_305), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_288), .ZN(n_0_0_306));
   OAI22_X1 i_0_0_402 (.A1(n_0_0_306), .A2(shift[0]), .B1(n_0_0_298), .B2(
      n_0_0_19), .ZN(n_0_125));
   AOI22_X1 i_0_0_403 (.A1(n_0_0_197), .A2(read_data2[18]), .B1(n_0_0_200), 
      .B2(n_0_51), .ZN(n_0_0_307));
   AOI22_X1 i_0_0_404 (.A1(n_0_0_196), .A2(n_0_21), .B1(read_data2[17]), 
      .B2(n_0_0_192), .ZN(n_0_0_308));
   NAND2_X1 i_0_0_405 (.A1(n_0_0_307), .A2(n_0_0_308), .ZN(n_0_0_309));
   OAI22_X1 i_0_0_406 (.A1(n_0_0_203), .A2(n_0_0_173), .B1(n_0_0_309), .B2(
      shift[4]), .ZN(n_0_0_310));
   INV_X1 i_0_0_407 (.A(n_0_0_310), .ZN(n_0_0_311));
   AOI22_X1 i_0_0_408 (.A1(n_0_0_311), .A2(n_0_0_172), .B1(n_0_0_256), .B2(
      n_0_0_244), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_409 (.A1(n_0_0_312), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_281), .ZN(n_0_0_313));
   AOI22_X1 i_0_0_410 (.A1(n_0_0_297), .A2(shift[1]), .B1(n_0_0_313), .B2(
      n_0_0_24), .ZN(n_0_0_314));
   OAI22_X1 i_0_0_411 (.A1(n_0_0_314), .A2(shift[0]), .B1(n_0_0_306), .B2(
      n_0_0_19), .ZN(n_0_126));
   AOI22_X1 i_0_0_412 (.A1(n_0_0_197), .A2(read_data2[19]), .B1(n_0_0_200), 
      .B2(n_0_52), .ZN(n_0_0_315));
   AOI22_X1 i_0_0_413 (.A1(n_0_0_196), .A2(n_0_22), .B1(read_data2[18]), 
      .B2(n_0_0_192), .ZN(n_0_0_316));
   NAND2_X1 i_0_0_414 (.A1(n_0_0_315), .A2(n_0_0_316), .ZN(n_0_0_317));
   OAI22_X1 i_0_0_415 (.A1(n_0_0_209), .A2(n_0_0_173), .B1(n_0_0_317), .B2(
      shift[4]), .ZN(n_0_0_318));
   NOR2_X1 i_0_0_416 (.A1(n_0_0_318), .A2(shift[5]), .ZN(n_0_0_319));
   AOI22_X1 i_0_0_417 (.A1(n_0_0_319), .A2(n_0_0_295), .B1(n_0_0_262), .B2(
      n_0_0_244), .ZN(n_0_0_320));
   OAI22_X1 i_0_0_418 (.A1(n_0_0_320), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_287), .ZN(n_0_0_321));
   AOI22_X1 i_0_0_419 (.A1(n_0_0_305), .A2(shift[1]), .B1(n_0_0_321), .B2(
      n_0_0_24), .ZN(n_0_0_322));
   OAI22_X1 i_0_0_420 (.A1(n_0_0_19), .A2(n_0_0_314), .B1(n_0_0_322), .B2(
      shift[0]), .ZN(n_0_127));
   AOI22_X1 i_0_0_421 (.A1(n_0_0_197), .A2(read_data2[20]), .B1(n_0_0_200), 
      .B2(n_0_53), .ZN(n_0_0_323));
   AOI22_X1 i_0_0_422 (.A1(n_0_0_196), .A2(n_0_23), .B1(read_data2[19]), 
      .B2(n_0_0_192), .ZN(n_0_0_324));
   NAND2_X1 i_0_0_423 (.A1(n_0_0_323), .A2(n_0_0_324), .ZN(n_0_0_325));
   OAI22_X1 i_0_0_424 (.A1(n_0_0_214), .A2(n_0_0_173), .B1(n_0_0_325), .B2(
      shift[4]), .ZN(n_0_0_326));
   INV_X1 i_0_0_425 (.A(n_0_0_326), .ZN(n_0_0_327));
   AOI22_X1 i_0_0_426 (.A1(n_0_0_327), .A2(n_0_0_172), .B1(n_0_0_268), .B2(
      n_0_0_244), .ZN(n_0_0_328));
   OAI22_X1 i_0_0_427 (.A1(n_0_0_328), .A2(shift[2]), .B1(n_0_0_296), .B2(
      n_0_0_23), .ZN(n_0_0_329));
   AOI22_X1 i_0_0_428 (.A1(n_0_0_329), .A2(n_0_0_24), .B1(n_0_0_313), .B2(
      shift[1]), .ZN(n_0_0_330));
   OAI22_X1 i_0_0_429 (.A1(shift[0]), .A2(n_0_0_330), .B1(n_0_0_322), .B2(
      n_0_0_19), .ZN(n_0_128));
   AOI22_X1 i_0_0_430 (.A1(n_0_0_197), .A2(read_data2[21]), .B1(n_0_0_200), 
      .B2(n_0_54), .ZN(n_0_0_331));
   AOI22_X1 i_0_0_431 (.A1(n_0_0_196), .A2(n_0_24), .B1(read_data2[20]), 
      .B2(n_0_0_192), .ZN(n_0_0_332));
   NAND2_X1 i_0_0_432 (.A1(n_0_0_331), .A2(n_0_0_332), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_433 (.A1(n_0_0_221), .A2(n_0_0_173), .B1(n_0_0_333), .B2(
      shift[4]), .ZN(n_0_0_334));
   INV_X1 i_0_0_434 (.A(n_0_0_334), .ZN(n_0_0_335));
   AOI22_X1 i_0_0_435 (.A1(n_0_0_335), .A2(n_0_0_172), .B1(n_0_0_274), .B2(
      n_0_0_244), .ZN(n_0_0_336));
   OAI22_X1 i_0_0_436 (.A1(n_0_0_304), .A2(n_0_0_23), .B1(n_0_0_336), .B2(
      shift[2]), .ZN(n_0_0_337));
   AOI22_X1 i_0_0_437 (.A1(n_0_0_337), .A2(n_0_0_24), .B1(n_0_0_321), .B2(
      shift[1]), .ZN(n_0_0_338));
   OAI22_X1 i_0_0_438 (.A1(n_0_0_338), .A2(shift[0]), .B1(n_0_0_330), .B2(
      n_0_0_19), .ZN(n_0_129));
   AOI22_X1 i_0_0_439 (.A1(n_0_0_197), .A2(read_data2[22]), .B1(n_0_0_200), 
      .B2(n_0_55), .ZN(n_0_0_339));
   AOI22_X1 i_0_0_440 (.A1(n_0_0_196), .A2(n_0_25), .B1(read_data2[21]), 
      .B2(n_0_0_192), .ZN(n_0_0_340));
   NAND2_X1 i_0_0_441 (.A1(n_0_0_339), .A2(n_0_0_340), .ZN(n_0_0_341));
   OAI22_X1 i_0_0_442 (.A1(n_0_0_228), .A2(n_0_0_173), .B1(n_0_0_341), .B2(
      shift[4]), .ZN(n_0_0_342));
   INV_X1 i_0_0_443 (.A(n_0_0_342), .ZN(n_0_0_343));
   AOI22_X1 i_0_0_444 (.A1(n_0_0_343), .A2(n_0_0_172), .B1(n_0_0_280), .B2(
      n_0_0_244), .ZN(n_0_0_344));
   OAI22_X1 i_0_0_445 (.A1(n_0_0_312), .A2(n_0_0_23), .B1(n_0_0_344), .B2(
      shift[2]), .ZN(n_0_0_345));
   AOI22_X1 i_0_0_446 (.A1(n_0_0_329), .A2(shift[1]), .B1(n_0_0_345), .B2(
      n_0_0_24), .ZN(n_0_0_346));
   OAI22_X1 i_0_0_447 (.A1(n_0_0_346), .A2(shift[0]), .B1(n_0_0_338), .B2(
      n_0_0_19), .ZN(n_0_130));
   AOI22_X1 i_0_0_448 (.A1(n_0_0_197), .A2(read_data2[23]), .B1(n_0_0_200), 
      .B2(n_0_56), .ZN(n_0_0_347));
   AOI22_X1 i_0_0_449 (.A1(n_0_0_196), .A2(n_0_26), .B1(read_data2[22]), 
      .B2(n_0_0_192), .ZN(n_0_0_348));
   NAND2_X1 i_0_0_450 (.A1(n_0_0_347), .A2(n_0_0_348), .ZN(n_0_0_349));
   OAI22_X1 i_0_0_451 (.A1(n_0_0_349), .A2(shift[4]), .B1(n_0_0_234), .B2(
      n_0_0_173), .ZN(n_0_0_350));
   INV_X1 i_0_0_452 (.A(n_0_0_350), .ZN(n_0_0_351));
   AOI22_X1 i_0_0_453 (.A1(n_0_0_351), .A2(n_0_0_172), .B1(n_0_0_286), .B2(
      n_0_0_244), .ZN(n_0_0_352));
   OAI22_X1 i_0_0_454 (.A1(n_0_0_352), .A2(shift[2]), .B1(n_0_0_320), .B2(
      n_0_0_23), .ZN(n_0_0_353));
   AOI22_X1 i_0_0_455 (.A1(n_0_0_337), .A2(shift[1]), .B1(n_0_0_353), .B2(
      n_0_0_24), .ZN(n_0_0_354));
   OAI22_X1 i_0_0_456 (.A1(n_0_0_346), .A2(n_0_0_19), .B1(n_0_0_354), .B2(
      shift[0]), .ZN(n_0_131));
   AOI22_X1 i_0_0_457 (.A1(n_0_0_196), .A2(n_0_27), .B1(n_0_0_200), .B2(n_0_57), 
      .ZN(n_0_0_355));
   AOI22_X1 i_0_0_458 (.A1(n_0_0_197), .A2(read_data2[24]), .B1(read_data2[23]), 
      .B2(n_0_0_192), .ZN(n_0_0_356));
   NAND2_X1 i_0_0_459 (.A1(n_0_0_355), .A2(n_0_0_356), .ZN(n_0_0_357));
   AOI22_X1 i_0_0_460 (.A1(n_0_0_357), .A2(n_0_0_173), .B1(n_0_0_241), .B2(
      shift[4]), .ZN(n_0_0_358));
   INV_X1 i_0_0_461 (.A(n_0_0_358), .ZN(n_0_0_359));
   AOI22_X1 i_0_0_462 (.A1(n_0_0_294), .A2(shift[3]), .B1(n_0_0_359), .B2(
      n_0_0_172), .ZN(n_0_0_360));
   OAI22_X1 i_0_0_463 (.A1(n_0_0_360), .A2(shift[2]), .B1(n_0_0_328), .B2(
      n_0_0_23), .ZN(n_0_0_361));
   AOI22_X1 i_0_0_464 (.A1(n_0_0_361), .A2(n_0_0_24), .B1(n_0_0_345), .B2(
      shift[1]), .ZN(n_0_0_362));
   OAI22_X1 i_0_0_465 (.A1(n_0_0_362), .A2(shift[0]), .B1(n_0_0_354), .B2(
      n_0_0_19), .ZN(n_0_132));
   INV_X1 i_0_0_466 (.A(n_0_0_243), .ZN(n_0_0_363));
   AOI22_X1 i_0_0_467 (.A1(n_0_0_197), .A2(read_data2[25]), .B1(n_0_0_200), 
      .B2(n_0_58), .ZN(n_0_0_364));
   AOI22_X1 i_0_0_468 (.A1(n_0_0_196), .A2(n_0_28), .B1(read_data2[24]), 
      .B2(n_0_0_192), .ZN(n_0_0_365));
   NAND2_X1 i_0_0_469 (.A1(n_0_0_364), .A2(n_0_0_365), .ZN(n_0_0_366));
   OAI22_X1 i_0_0_470 (.A1(n_0_0_250), .A2(n_0_0_173), .B1(n_0_0_366), .B2(
      shift[4]), .ZN(n_0_0_367));
   INV_X1 i_0_0_471 (.A(n_0_0_367), .ZN(n_0_0_368));
   AOI22_X1 i_0_0_472 (.A1(n_0_0_303), .A2(n_0_0_363), .B1(n_0_0_368), .B2(
      n_0_0_172), .ZN(n_0_0_369));
   OAI22_X1 i_0_0_473 (.A1(n_0_0_369), .A2(shift[2]), .B1(n_0_0_336), .B2(
      n_0_0_23), .ZN(n_0_0_370));
   AOI22_X1 i_0_0_474 (.A1(n_0_0_370), .A2(n_0_0_24), .B1(n_0_0_353), .B2(
      shift[1]), .ZN(n_0_0_371));
   OAI22_X1 i_0_0_475 (.A1(n_0_0_362), .A2(n_0_0_19), .B1(n_0_0_371), .B2(
      shift[0]), .ZN(n_0_133));
   AOI22_X1 i_0_0_476 (.A1(n_0_0_196), .A2(n_0_29), .B1(n_0_0_200), .B2(n_0_59), 
      .ZN(n_0_0_372));
   AOI22_X1 i_0_0_477 (.A1(n_0_0_197), .A2(read_data2[26]), .B1(read_data2[25]), 
      .B2(n_0_0_192), .ZN(n_0_0_373));
   NAND2_X1 i_0_0_478 (.A1(n_0_0_372), .A2(n_0_0_373), .ZN(n_0_0_374));
   OAI22_X1 i_0_0_479 (.A1(n_0_0_374), .A2(shift[4]), .B1(n_0_0_256), .B2(
      n_0_0_173), .ZN(n_0_0_375));
   INV_X1 i_0_0_480 (.A(n_0_0_375), .ZN(n_0_0_376));
   AOI22_X1 i_0_0_481 (.A1(n_0_0_311), .A2(n_0_0_363), .B1(n_0_0_376), .B2(
      n_0_0_172), .ZN(n_0_0_377));
   OAI22_X1 i_0_0_482 (.A1(n_0_0_377), .A2(shift[2]), .B1(n_0_0_344), .B2(
      n_0_0_23), .ZN(n_0_0_378));
   AOI22_X1 i_0_0_483 (.A1(n_0_0_361), .A2(shift[1]), .B1(n_0_0_378), .B2(
      n_0_0_24), .ZN(n_0_0_379));
   OAI22_X1 i_0_0_484 (.A1(n_0_0_379), .A2(shift[0]), .B1(n_0_0_371), .B2(
      n_0_0_19), .ZN(n_0_134));
   INV_X1 i_0_0_485 (.A(n_0_0_262), .ZN(n_0_0_380));
   AOI22_X1 i_0_0_486 (.A1(n_0_0_196), .A2(n_0_30), .B1(n_0_0_200), .B2(n_0_60), 
      .ZN(n_0_0_381));
   AOI22_X1 i_0_0_487 (.A1(n_0_0_197), .A2(read_data2[27]), .B1(read_data2[26]), 
      .B2(n_0_0_192), .ZN(n_0_0_382));
   AND2_X1 i_0_0_488 (.A1(n_0_0_381), .A2(n_0_0_382), .ZN(n_0_0_383));
   AOI22_X1 i_0_0_489 (.A1(n_0_0_380), .A2(shift[4]), .B1(n_0_0_383), .B2(
      n_0_0_173), .ZN(n_0_0_384));
   AOI22_X1 i_0_0_490 (.A1(n_0_0_319), .A2(shift[3]), .B1(n_0_0_384), .B2(
      n_0_0_172), .ZN(n_0_0_385));
   OAI22_X1 i_0_0_491 (.A1(n_0_0_385), .A2(shift[2]), .B1(n_0_0_352), .B2(
      n_0_0_23), .ZN(n_0_0_386));
   AOI22_X1 i_0_0_492 (.A1(n_0_0_370), .A2(shift[1]), .B1(n_0_0_386), .B2(
      n_0_0_24), .ZN(n_0_0_387));
   OAI22_X1 i_0_0_493 (.A1(n_0_0_387), .A2(shift[0]), .B1(n_0_0_379), .B2(
      n_0_0_19), .ZN(n_0_135));
   INV_X1 i_0_0_494 (.A(n_0_0_268), .ZN(n_0_0_388));
   NAND2_X1 i_0_0_495 (.A1(n_0_0_33), .A2(shift[4]), .ZN(n_0_0_389));
   AOI22_X1 i_0_0_496 (.A1(n_0_0_197), .A2(read_data2[28]), .B1(n_0_0_200), 
      .B2(n_0_61), .ZN(n_0_0_390));
   AOI22_X1 i_0_0_497 (.A1(n_0_0_196), .A2(n_0_31), .B1(read_data2[27]), 
      .B2(n_0_0_192), .ZN(n_0_0_391));
   AND2_X1 i_0_0_498 (.A1(n_0_0_390), .A2(n_0_0_391), .ZN(n_0_0_392));
   NAND2_X1 i_0_0_499 (.A1(n_0_0_173), .A2(n_0_0_33), .ZN(n_0_0_393));
   OAI22_X1 i_0_0_500 (.A1(n_0_0_388), .A2(n_0_0_389), .B1(n_0_0_392), .B2(
      n_0_0_393), .ZN(n_0_0_394));
   AOI22_X1 i_0_0_501 (.A1(n_0_0_394), .A2(n_0_0_295), .B1(n_0_0_327), .B2(
      n_0_0_363), .ZN(n_0_0_395));
   OAI22_X1 i_0_0_502 (.A1(n_0_0_395), .A2(shift[2]), .B1(n_0_0_360), .B2(
      n_0_0_23), .ZN(n_0_0_396));
   AOI22_X1 i_0_0_503 (.A1(n_0_0_396), .A2(n_0_0_24), .B1(n_0_0_378), .B2(
      shift[1]), .ZN(n_0_0_397));
   OAI22_X1 i_0_0_504 (.A1(n_0_0_387), .A2(n_0_0_19), .B1(n_0_0_397), .B2(
      shift[0]), .ZN(n_0_136));
   INV_X1 i_0_0_505 (.A(n_0_0_274), .ZN(n_0_0_398));
   AOI22_X1 i_0_0_506 (.A1(n_0_0_197), .A2(read_data2[29]), .B1(n_0_0_200), 
      .B2(n_0_62), .ZN(n_0_0_399));
   AOI22_X1 i_0_0_507 (.A1(n_0_0_196), .A2(n_0_32), .B1(read_data2[28]), 
      .B2(n_0_0_192), .ZN(n_0_0_400));
   AND2_X1 i_0_0_508 (.A1(n_0_0_399), .A2(n_0_0_400), .ZN(n_0_0_401));
   OAI22_X1 i_0_0_509 (.A1(n_0_0_398), .A2(n_0_0_173), .B1(n_0_0_401), .B2(
      shift[4]), .ZN(n_0_0_402));
   AOI22_X1 i_0_0_510 (.A1(n_0_0_335), .A2(n_0_0_363), .B1(n_0_0_402), .B2(
      n_0_0_172), .ZN(n_0_0_403));
   OAI22_X1 i_0_0_511 (.A1(n_0_0_369), .A2(n_0_0_23), .B1(n_0_0_403), .B2(
      shift[2]), .ZN(n_0_0_404));
   AOI22_X1 i_0_0_512 (.A1(n_0_0_404), .A2(n_0_0_24), .B1(n_0_0_386), .B2(
      shift[1]), .ZN(n_0_0_405));
   OAI22_X1 i_0_0_513 (.A1(n_0_0_405), .A2(shift[0]), .B1(n_0_0_397), .B2(
      n_0_0_19), .ZN(n_0_137));
   INV_X1 i_0_0_514 (.A(n_0_0_280), .ZN(n_0_0_406));
   AOI22_X1 i_0_0_515 (.A1(n_0_0_196), .A2(n_0_33), .B1(n_0_0_200), .B2(n_0_63), 
      .ZN(n_0_0_407));
   AOI22_X1 i_0_0_516 (.A1(n_0_0_197), .A2(read_data2[30]), .B1(read_data2[29]), 
      .B2(n_0_0_192), .ZN(n_0_0_408));
   AND2_X1 i_0_0_517 (.A1(n_0_0_407), .A2(n_0_0_408), .ZN(n_0_0_409));
   OAI22_X1 i_0_0_518 (.A1(n_0_0_406), .A2(n_0_0_173), .B1(n_0_0_409), .B2(
      shift[4]), .ZN(n_0_0_410));
   AOI22_X1 i_0_0_519 (.A1(n_0_0_343), .A2(n_0_0_363), .B1(n_0_0_410), .B2(
      n_0_0_172), .ZN(n_0_0_411));
   OAI22_X1 i_0_0_520 (.A1(n_0_0_377), .A2(n_0_0_23), .B1(n_0_0_411), .B2(
      shift[2]), .ZN(n_0_0_412));
   AOI22_X1 i_0_0_521 (.A1(n_0_0_396), .A2(shift[1]), .B1(n_0_0_412), .B2(
      n_0_0_24), .ZN(n_0_0_413));
   OAI22_X1 i_0_0_522 (.A1(n_0_0_405), .A2(n_0_0_19), .B1(n_0_0_413), .B2(
      shift[0]), .ZN(n_0_138));
   AOI22_X1 i_0_0_523 (.A1(n_0_0_196), .A2(n_0_34), .B1(n_0_0_197), .B2(
      read_data2[31]), .ZN(n_0_0_414));
   AOI22_X1 i_0_0_524 (.A1(n_0_0_200), .A2(n_0_64), .B1(read_data2[30]), 
      .B2(n_0_0_192), .ZN(n_0_0_415));
   AND2_X1 i_0_0_525 (.A1(n_0_0_414), .A2(n_0_0_415), .ZN(n_0_0_416));
   INV_X1 i_0_0_526 (.A(n_0_0_286), .ZN(n_0_0_417));
   OAI22_X1 i_0_0_527 (.A1(n_0_0_416), .A2(n_0_0_393), .B1(n_0_0_417), .B2(
      n_0_0_389), .ZN(n_0_0_418));
   AOI22_X1 i_0_0_528 (.A1(n_0_0_418), .A2(n_0_0_295), .B1(n_0_0_351), .B2(
      n_0_0_363), .ZN(n_0_0_419));
   OAI22_X1 i_0_0_529 (.A1(n_0_0_385), .A2(n_0_0_23), .B1(n_0_0_419), .B2(
      shift[2]), .ZN(n_0_0_420));
   AOI22_X1 i_0_0_530 (.A1(n_0_0_404), .A2(shift[1]), .B1(n_0_0_420), .B2(
      n_0_0_24), .ZN(n_0_0_421));
   OAI22_X1 i_0_0_531 (.A1(n_0_0_421), .A2(shift[0]), .B1(n_0_0_413), .B2(
      n_0_0_19), .ZN(n_0_139));
   AOI22_X1 i_0_0_532 (.A1(n_0_0_200), .A2(n_0_65), .B1(read_data2[31]), 
      .B2(n_0_0_192), .ZN(n_0_0_422));
   NAND2_X1 i_0_0_533 (.A1(n_0_0_414), .A2(n_0_0_422), .ZN(n_0_107));
   AND2_X1 i_0_0_534 (.A1(n_0_107), .A2(n_0_0_33), .ZN(n_0_0_423));
   INV_X1 i_0_0_535 (.A(n_0_0_423), .ZN(n_0_0_424));
   NOR2_X1 i_0_0_536 (.A1(n_0_0_424), .A2(shift[4]), .ZN(n_0_0_425));
   INV_X1 i_0_0_537 (.A(n_0_0_389), .ZN(n_0_0_426));
   AOI21_X1 i_0_0_538 (.A(n_0_0_425), .B1(n_0_0_292), .B2(n_0_0_426), .ZN(
      n_0_0_427));
   NAND2_X1 i_0_0_539 (.A1(n_0_0_173), .A2(shift[5]), .ZN(n_0_0_428));
   OAI21_X1 i_0_0_540 (.A(n_0_0_427), .B1(n_0_0_171), .B2(n_0_0_428), .ZN(
      n_0_0_429));
   AOI22_X1 i_0_0_541 (.A1(n_0_0_429), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_359), .ZN(n_0_0_430));
   OAI22_X1 i_0_0_542 (.A1(n_0_0_430), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_395), .ZN(n_0_0_431));
   AOI22_X1 i_0_0_543 (.A1(n_0_0_431), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_412), .ZN(n_0_0_432));
   OAI22_X1 i_0_0_544 (.A1(n_0_0_432), .A2(shift[0]), .B1(n_0_0_421), .B2(
      n_0_0_19), .ZN(n_0_140));
   INV_X1 i_0_0_545 (.A(n_0_0_425), .ZN(n_0_0_433));
   INV_X1 i_0_0_546 (.A(n_0_0_301), .ZN(n_0_0_434));
   OAI221_X1 i_0_0_547 (.A(n_0_0_433), .B1(n_0_0_434), .B2(n_0_0_389), .C1(
      n_0_0_198), .C2(n_0_0_428), .ZN(n_0_0_435));
   AOI22_X1 i_0_0_548 (.A1(n_0_0_435), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_368), .ZN(n_0_0_436));
   OAI22_X1 i_0_0_549 (.A1(n_0_0_436), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_403), .ZN(n_0_0_437));
   AOI22_X1 i_0_0_550 (.A1(n_0_0_437), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_420), .ZN(n_0_0_438));
   OAI22_X1 i_0_0_551 (.A1(n_0_0_438), .A2(shift[0]), .B1(n_0_0_19), .B2(
      n_0_0_432), .ZN(n_0_141));
   INV_X1 i_0_0_552 (.A(n_0_0_309), .ZN(n_0_0_439));
   OAI221_X1 i_0_0_553 (.A(n_0_0_433), .B1(n_0_0_225), .B2(n_0_0_428), .C1(
      n_0_0_439), .C2(n_0_0_389), .ZN(n_0_0_440));
   AOI22_X1 i_0_0_554 (.A1(n_0_0_440), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_376), .ZN(n_0_0_441));
   OAI22_X1 i_0_0_555 (.A1(n_0_0_441), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_411), .ZN(n_0_0_442));
   AOI22_X1 i_0_0_556 (.A1(n_0_0_442), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_431), .ZN(n_0_0_443));
   OAI22_X1 i_0_0_557 (.A1(n_0_0_443), .A2(shift[0]), .B1(n_0_0_438), .B2(
      n_0_0_19), .ZN(n_0_142));
   INV_X1 i_0_0_558 (.A(n_0_0_317), .ZN(n_0_0_444));
   OAI221_X1 i_0_0_559 (.A(n_0_0_433), .B1(n_0_0_236), .B2(n_0_0_428), .C1(
      n_0_0_444), .C2(n_0_0_389), .ZN(n_0_0_445));
   AOI22_X1 i_0_0_560 (.A1(n_0_0_445), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_384), .ZN(n_0_0_446));
   OAI22_X1 i_0_0_561 (.A1(n_0_0_446), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_419), .ZN(n_0_0_447));
   AOI22_X1 i_0_0_562 (.A1(n_0_0_437), .A2(shift[1]), .B1(n_0_0_447), .B2(
      n_0_0_24), .ZN(n_0_0_448));
   OAI22_X1 i_0_0_563 (.A1(n_0_0_448), .A2(shift[0]), .B1(n_0_0_443), .B2(
      n_0_0_19), .ZN(n_0_143));
   INV_X1 i_0_0_564 (.A(n_0_0_325), .ZN(n_0_0_449));
   OAI221_X1 i_0_0_565 (.A(n_0_0_433), .B1(n_0_0_215), .B2(n_0_0_428), .C1(
      n_0_0_449), .C2(n_0_0_389), .ZN(n_0_0_450));
   AOI22_X1 i_0_0_566 (.A1(n_0_0_450), .A2(n_0_0_295), .B1(shift[3]), .B2(
      n_0_0_394), .ZN(n_0_0_451));
   OAI22_X1 i_0_0_567 (.A1(n_0_0_451), .A2(shift[2]), .B1(n_0_0_23), .B2(
      n_0_0_430), .ZN(n_0_0_452));
   AOI22_X1 i_0_0_568 (.A1(n_0_0_452), .A2(n_0_0_24), .B1(n_0_0_442), .B2(
      shift[1]), .ZN(n_0_0_453));
   OAI22_X1 i_0_0_569 (.A1(n_0_0_448), .A2(n_0_0_19), .B1(n_0_0_453), .B2(
      shift[0]), .ZN(n_0_144));
   INV_X1 i_0_0_570 (.A(n_0_0_333), .ZN(n_0_0_454));
   OAI221_X1 i_0_0_571 (.A(n_0_0_433), .B1(n_0_0_222), .B2(n_0_0_428), .C1(
      n_0_0_454), .C2(n_0_0_389), .ZN(n_0_0_455));
   AOI22_X1 i_0_0_572 (.A1(n_0_0_455), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_402), .ZN(n_0_0_456));
   OAI22_X1 i_0_0_573 (.A1(n_0_0_436), .A2(n_0_0_23), .B1(n_0_0_456), .B2(
      shift[2]), .ZN(n_0_0_457));
   AOI22_X1 i_0_0_574 (.A1(n_0_0_457), .A2(n_0_0_24), .B1(n_0_0_447), .B2(
      shift[1]), .ZN(n_0_0_458));
   OAI22_X1 i_0_0_575 (.A1(n_0_0_458), .A2(shift[0]), .B1(n_0_0_453), .B2(
      n_0_0_19), .ZN(n_0_145));
   INV_X1 i_0_0_576 (.A(n_0_0_341), .ZN(n_0_0_459));
   OAI221_X1 i_0_0_577 (.A(n_0_0_433), .B1(n_0_0_229), .B2(n_0_0_428), .C1(
      n_0_0_459), .C2(n_0_0_389), .ZN(n_0_0_460));
   AOI22_X1 i_0_0_578 (.A1(n_0_0_460), .A2(n_0_0_295), .B1(n_0_0_363), .B2(
      n_0_0_410), .ZN(n_0_0_461));
   OAI22_X1 i_0_0_579 (.A1(n_0_0_461), .A2(shift[2]), .B1(n_0_0_441), .B2(
      n_0_0_23), .ZN(n_0_0_462));
   AOI22_X1 i_0_0_580 (.A1(n_0_0_462), .A2(n_0_0_24), .B1(n_0_0_452), .B2(
      shift[1]), .ZN(n_0_0_463));
   OAI22_X1 i_0_0_581 (.A1(n_0_0_463), .A2(shift[0]), .B1(n_0_0_458), .B2(
      n_0_0_19), .ZN(n_0_146));
   INV_X1 i_0_0_582 (.A(n_0_0_349), .ZN(n_0_0_464));
   OAI221_X1 i_0_0_583 (.A(n_0_0_433), .B1(n_0_0_464), .B2(n_0_0_389), .C1(
      n_0_0_235), .C2(n_0_0_428), .ZN(n_0_0_465));
   AOI22_X1 i_0_0_584 (.A1(n_0_0_465), .A2(n_0_0_295), .B1(shift[3]), .B2(
      n_0_0_418), .ZN(n_0_0_466));
   OAI22_X1 i_0_0_585 (.A1(n_0_0_466), .A2(shift[2]), .B1(n_0_0_446), .B2(
      n_0_0_23), .ZN(n_0_0_467));
   AOI22_X1 i_0_0_586 (.A1(n_0_0_457), .A2(shift[1]), .B1(n_0_0_467), .B2(
      n_0_0_24), .ZN(n_0_0_468));
   OAI22_X1 i_0_0_587 (.A1(n_0_0_468), .A2(shift[0]), .B1(n_0_0_463), .B2(
      n_0_0_19), .ZN(n_0_147));
   INV_X1 i_0_0_588 (.A(n_0_0_241), .ZN(n_0_0_469));
   INV_X1 i_0_0_589 (.A(n_0_0_357), .ZN(n_0_0_470));
   OAI221_X1 i_0_0_590 (.A(n_0_0_433), .B1(n_0_0_469), .B2(n_0_0_428), .C1(
      n_0_0_470), .C2(n_0_0_389), .ZN(n_0_0_471));
   AOI22_X1 i_0_0_591 (.A1(n_0_0_471), .A2(n_0_0_295), .B1(n_0_0_429), .B2(
      shift[3]), .ZN(n_0_0_472));
   OAI22_X1 i_0_0_592 (.A1(n_0_0_451), .A2(n_0_0_23), .B1(n_0_0_472), .B2(
      shift[2]), .ZN(n_0_0_473));
   AOI22_X1 i_0_0_593 (.A1(n_0_0_462), .A2(shift[1]), .B1(n_0_0_473), .B2(
      n_0_0_24), .ZN(n_0_0_474));
   OAI22_X1 i_0_0_594 (.A1(n_0_0_468), .A2(n_0_0_19), .B1(n_0_0_474), .B2(
      shift[0]), .ZN(n_0_148));
   INV_X1 i_0_0_595 (.A(n_0_0_366), .ZN(n_0_0_475));
   INV_X1 i_0_0_596 (.A(n_0_0_250), .ZN(n_0_0_476));
   OAI221_X1 i_0_0_597 (.A(n_0_0_433), .B1(n_0_0_475), .B2(n_0_0_389), .C1(
      n_0_0_476), .C2(n_0_0_428), .ZN(n_0_0_477));
   OAI22_X1 i_0_0_598 (.A1(n_0_0_477), .A2(shift[3]), .B1(n_0_0_435), .B2(
      n_0_0_295), .ZN(n_0_0_478));
   AOI22_X1 i_0_0_599 (.A1(n_0_0_478), .A2(n_0_0_23), .B1(n_0_0_456), .B2(
      shift[2]), .ZN(n_0_0_479));
   AOI22_X1 i_0_0_600 (.A1(n_0_0_479), .A2(n_0_0_24), .B1(n_0_0_467), .B2(
      shift[1]), .ZN(n_0_0_480));
   OAI22_X1 i_0_0_601 (.A1(n_0_0_480), .A2(shift[0]), .B1(n_0_0_474), .B2(
      n_0_0_19), .ZN(n_0_149));
   INV_X1 i_0_0_602 (.A(n_0_0_256), .ZN(n_0_0_481));
   INV_X1 i_0_0_603 (.A(n_0_0_374), .ZN(n_0_0_482));
   OAI221_X1 i_0_0_604 (.A(n_0_0_433), .B1(n_0_0_481), .B2(n_0_0_428), .C1(
      n_0_0_482), .C2(n_0_0_389), .ZN(n_0_0_483));
   AOI22_X1 i_0_0_605 (.A1(n_0_0_440), .A2(shift[3]), .B1(n_0_0_483), .B2(
      n_0_0_295), .ZN(n_0_0_484));
   OAI22_X1 i_0_0_606 (.A1(n_0_0_484), .A2(shift[2]), .B1(n_0_0_461), .B2(
      n_0_0_23), .ZN(n_0_0_485));
   AOI22_X1 i_0_0_607 (.A1(n_0_0_485), .A2(n_0_0_24), .B1(n_0_0_473), .B2(
      shift[1]), .ZN(n_0_0_486));
   OAI22_X1 i_0_0_608 (.A1(n_0_0_480), .A2(n_0_0_19), .B1(n_0_0_486), .B2(
      shift[0]), .ZN(n_0_150));
   OAI221_X1 i_0_0_609 (.A(n_0_0_433), .B1(n_0_0_383), .B2(n_0_0_389), .C1(
      n_0_0_380), .C2(n_0_0_428), .ZN(n_0_0_487));
   OAI22_X1 i_0_0_610 (.A1(n_0_0_445), .A2(n_0_0_295), .B1(n_0_0_487), .B2(
      shift[3]), .ZN(n_0_0_488));
   OAI22_X1 i_0_0_611 (.A1(n_0_0_488), .A2(shift[2]), .B1(n_0_0_466), .B2(
      n_0_0_23), .ZN(n_0_0_489));
   AOI22_X1 i_0_0_612 (.A1(n_0_0_479), .A2(shift[1]), .B1(n_0_0_489), .B2(
      n_0_0_24), .ZN(n_0_0_490));
   OAI22_X1 i_0_0_613 (.A1(n_0_0_490), .A2(shift[0]), .B1(n_0_0_486), .B2(
      n_0_0_19), .ZN(n_0_151));
   AOI21_X1 i_0_0_614 (.A(n_0_0_423), .B1(shift[5]), .B2(n_0_0_268), .ZN(
      n_0_0_491));
   OAI22_X1 i_0_0_615 (.A1(n_0_0_491), .A2(shift[4]), .B1(n_0_0_389), .B2(
      n_0_0_392), .ZN(n_0_0_492));
   AOI22_X1 i_0_0_616 (.A1(n_0_0_450), .A2(shift[3]), .B1(n_0_0_492), .B2(
      n_0_0_295), .ZN(n_0_0_493));
   OAI22_X1 i_0_0_617 (.A1(n_0_0_493), .A2(shift[2]), .B1(n_0_0_472), .B2(
      n_0_0_23), .ZN(n_0_0_494));
   AOI22_X1 i_0_0_618 (.A1(n_0_0_485), .A2(shift[1]), .B1(n_0_0_494), .B2(
      n_0_0_24), .ZN(n_0_0_495));
   OAI22_X1 i_0_0_619 (.A1(n_0_0_490), .A2(n_0_0_19), .B1(n_0_0_495), .B2(
      shift[0]), .ZN(n_0_152));
   OAI221_X1 i_0_0_620 (.A(n_0_0_433), .B1(n_0_0_398), .B2(n_0_0_428), .C1(
      n_0_0_389), .C2(n_0_0_401), .ZN(n_0_0_496));
   AOI22_X1 i_0_0_621 (.A1(n_0_0_455), .A2(shift[3]), .B1(n_0_0_496), .B2(
      n_0_0_295), .ZN(n_0_0_497));
   OAI22_X1 i_0_0_622 (.A1(n_0_0_497), .A2(shift[2]), .B1(n_0_0_478), .B2(
      n_0_0_23), .ZN(n_0_0_498));
   AOI22_X1 i_0_0_623 (.A1(n_0_0_498), .A2(n_0_0_24), .B1(n_0_0_489), .B2(
      shift[1]), .ZN(n_0_0_499));
   OAI22_X1 i_0_0_624 (.A1(n_0_0_499), .A2(shift[0]), .B1(n_0_0_495), .B2(
      n_0_0_19), .ZN(n_0_153));
   OAI221_X1 i_0_0_625 (.A(n_0_0_433), .B1(n_0_0_406), .B2(n_0_0_428), .C1(
      n_0_0_389), .C2(n_0_0_409), .ZN(n_0_0_500));
   AOI22_X1 i_0_0_626 (.A1(n_0_0_460), .A2(shift[3]), .B1(n_0_0_500), .B2(
      n_0_0_295), .ZN(n_0_0_501));
   OAI22_X1 i_0_0_627 (.A1(n_0_0_484), .A2(n_0_0_23), .B1(n_0_0_501), .B2(
      shift[2]), .ZN(n_0_0_502));
   AOI22_X1 i_0_0_628 (.A1(n_0_0_502), .A2(n_0_0_24), .B1(n_0_0_494), .B2(
      shift[1]), .ZN(n_0_0_503));
   OAI22_X1 i_0_0_629 (.A1(n_0_0_499), .A2(n_0_0_19), .B1(n_0_0_503), .B2(
      shift[0]), .ZN(n_0_154));
   OAI221_X1 i_0_0_630 (.A(n_0_0_433), .B1(n_0_0_417), .B2(n_0_0_428), .C1(
      n_0_0_389), .C2(n_0_0_416), .ZN(n_0_0_504));
   AOI22_X1 i_0_0_631 (.A1(n_0_0_465), .A2(shift[3]), .B1(n_0_0_504), .B2(
      n_0_0_295), .ZN(n_0_0_505));
   OAI22_X1 i_0_0_632 (.A1(n_0_0_505), .A2(shift[2]), .B1(n_0_0_488), .B2(
      n_0_0_23), .ZN(n_0_0_506));
   AOI22_X1 i_0_0_633 (.A1(n_0_0_498), .A2(shift[1]), .B1(n_0_0_506), .B2(
      n_0_0_24), .ZN(n_0_0_507));
   OAI22_X1 i_0_0_634 (.A1(n_0_0_507), .A2(shift[0]), .B1(n_0_0_503), .B2(
      n_0_0_19), .ZN(n_0_155));
   NOR2_X1 i_0_0_635 (.A1(n_0_0_423), .A2(shift[3]), .ZN(n_0_0_508));
   INV_X1 i_0_0_636 (.A(n_0_0_508), .ZN(n_0_0_509));
   NOR2_X1 i_0_0_637 (.A1(n_0_0_293), .A2(n_0_0_33), .ZN(n_0_0_510));
   OAI22_X1 i_0_0_638 (.A1(n_0_0_471), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_510), .ZN(n_0_0_511));
   OAI22_X1 i_0_0_639 (.A1(n_0_0_511), .A2(shift[2]), .B1(n_0_0_493), .B2(
      n_0_0_23), .ZN(n_0_0_512));
   AOI22_X1 i_0_0_640 (.A1(n_0_0_502), .A2(shift[1]), .B1(n_0_0_512), .B2(
      n_0_0_24), .ZN(n_0_0_513));
   OAI22_X1 i_0_0_641 (.A1(n_0_0_507), .A2(n_0_0_19), .B1(n_0_0_513), .B2(
      shift[0]), .ZN(n_0_156));
   NOR2_X1 i_0_0_642 (.A1(n_0_0_302), .A2(n_0_0_33), .ZN(n_0_0_514));
   OAI22_X1 i_0_0_643 (.A1(n_0_0_477), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_514), .ZN(n_0_0_515));
   OAI22_X1 i_0_0_644 (.A1(n_0_0_497), .A2(n_0_0_23), .B1(n_0_0_515), .B2(
      shift[2]), .ZN(n_0_0_516));
   AOI22_X1 i_0_0_645 (.A1(shift[1]), .A2(n_0_0_506), .B1(n_0_0_516), .B2(
      n_0_0_24), .ZN(n_0_0_517));
   OAI22_X1 i_0_0_646 (.A1(n_0_0_517), .A2(shift[0]), .B1(n_0_0_513), .B2(
      n_0_0_19), .ZN(n_0_157));
   NOR2_X1 i_0_0_647 (.A1(n_0_0_310), .A2(n_0_0_33), .ZN(n_0_0_518));
   OAI22_X1 i_0_0_648 (.A1(n_0_0_483), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_518), .ZN(n_0_0_519));
   OAI22_X1 i_0_0_649 (.A1(n_0_0_501), .A2(n_0_0_23), .B1(n_0_0_519), .B2(
      shift[2]), .ZN(n_0_0_520));
   AOI22_X1 i_0_0_650 (.A1(n_0_0_520), .A2(n_0_0_24), .B1(n_0_0_512), .B2(
      shift[1]), .ZN(n_0_0_521));
   OAI22_X1 i_0_0_651 (.A1(n_0_0_517), .A2(n_0_0_19), .B1(n_0_0_521), .B2(
      shift[0]), .ZN(n_0_158));
   NOR2_X1 i_0_0_652 (.A1(n_0_0_318), .A2(n_0_0_33), .ZN(n_0_0_522));
   OAI22_X1 i_0_0_653 (.A1(n_0_0_487), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_522), .ZN(n_0_0_523));
   OAI22_X1 i_0_0_654 (.A1(n_0_0_505), .A2(n_0_0_23), .B1(n_0_0_523), .B2(
      shift[2]), .ZN(n_0_0_524));
   AOI22_X1 i_0_0_655 (.A1(n_0_0_516), .A2(shift[1]), .B1(n_0_0_524), .B2(
      n_0_0_24), .ZN(n_0_0_525));
   OAI22_X1 i_0_0_656 (.A1(n_0_0_525), .A2(shift[0]), .B1(n_0_0_521), .B2(
      n_0_0_19), .ZN(n_0_159));
   NOR2_X1 i_0_0_657 (.A1(n_0_0_326), .A2(n_0_0_33), .ZN(n_0_0_526));
   OAI22_X1 i_0_0_658 (.A1(n_0_0_492), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_526), .ZN(n_0_0_527));
   OAI22_X1 i_0_0_659 (.A1(n_0_0_511), .A2(n_0_0_23), .B1(n_0_0_527), .B2(
      shift[2]), .ZN(n_0_0_528));
   AOI22_X1 i_0_0_660 (.A1(n_0_0_520), .A2(shift[1]), .B1(n_0_0_528), .B2(
      n_0_0_24), .ZN(n_0_0_529));
   OAI22_X1 i_0_0_661 (.A1(n_0_0_525), .A2(n_0_0_19), .B1(n_0_0_529), .B2(
      shift[0]), .ZN(n_0_160));
   NOR2_X1 i_0_0_662 (.A1(n_0_0_334), .A2(n_0_0_33), .ZN(n_0_0_530));
   OAI22_X1 i_0_0_663 (.A1(n_0_0_496), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_530), .ZN(n_0_0_531));
   AOI22_X1 i_0_0_664 (.A1(n_0_0_515), .A2(shift[2]), .B1(n_0_0_531), .B2(
      n_0_0_23), .ZN(n_0_0_532));
   AOI22_X1 i_0_0_665 (.A1(n_0_0_524), .A2(shift[1]), .B1(n_0_0_532), .B2(
      n_0_0_24), .ZN(n_0_0_533));
   OAI22_X1 i_0_0_666 (.A1(n_0_0_533), .A2(shift[0]), .B1(n_0_0_529), .B2(
      n_0_0_19), .ZN(n_0_161));
   NOR2_X1 i_0_0_667 (.A1(n_0_0_342), .A2(n_0_0_33), .ZN(n_0_0_534));
   OAI22_X1 i_0_0_668 (.A1(n_0_0_500), .A2(n_0_0_295), .B1(n_0_0_509), .B2(
      n_0_0_534), .ZN(n_0_0_535));
   OAI22_X1 i_0_0_669 (.A1(n_0_0_519), .A2(n_0_0_23), .B1(n_0_0_535), .B2(
      shift[2]), .ZN(n_0_0_536));
   AOI22_X1 i_0_0_670 (.A1(n_0_0_536), .A2(n_0_0_24), .B1(n_0_0_528), .B2(
      shift[1]), .ZN(n_0_0_537));
   OAI22_X1 i_0_0_671 (.A1(n_0_0_533), .A2(n_0_0_19), .B1(n_0_0_537), .B2(
      shift[0]), .ZN(n_0_162));
   OAI21_X1 i_0_0_672 (.A(n_0_0_508), .B1(n_0_0_33), .B2(n_0_0_350), .ZN(
      n_0_0_538));
   OAI21_X1 i_0_0_673 (.A(n_0_0_538), .B1(n_0_0_504), .B2(n_0_0_295), .ZN(
      n_0_0_539));
   OAI22_X1 i_0_0_674 (.A1(n_0_0_523), .A2(n_0_0_23), .B1(n_0_0_539), .B2(
      shift[2]), .ZN(n_0_0_540));
   OAI22_X1 i_0_0_675 (.A1(n_0_0_532), .A2(n_0_0_24), .B1(n_0_0_540), .B2(
      shift[1]), .ZN(n_0_0_541));
   OAI22_X1 i_0_0_676 (.A1(n_0_0_541), .A2(shift[0]), .B1(n_0_0_537), .B2(
      n_0_0_19), .ZN(n_0_163));
   NOR2_X1 i_0_0_677 (.A1(n_0_0_358), .A2(n_0_0_33), .ZN(n_0_0_542));
   NAND2_X1 i_0_0_678 (.A1(n_0_0_424), .A2(shift[3]), .ZN(n_0_0_543));
   OAI22_X1 i_0_0_679 (.A1(n_0_0_542), .A2(n_0_0_509), .B1(n_0_0_510), .B2(
      n_0_0_543), .ZN(n_0_0_544));
   OAI22_X1 i_0_0_680 (.A1(n_0_0_527), .A2(n_0_0_23), .B1(shift[2]), .B2(
      n_0_0_544), .ZN(n_0_0_545));
   AOI22_X1 i_0_0_681 (.A1(n_0_0_536), .A2(shift[1]), .B1(n_0_0_24), .B2(
      n_0_0_545), .ZN(n_0_0_546));
   OAI22_X1 i_0_0_682 (.A1(n_0_0_541), .A2(n_0_0_19), .B1(n_0_0_546), .B2(
      shift[0]), .ZN(n_0_164));
   NOR2_X1 i_0_0_683 (.A1(n_0_0_367), .A2(n_0_0_33), .ZN(n_0_0_547));
   OAI22_X1 i_0_0_684 (.A1(n_0_0_547), .A2(n_0_0_509), .B1(n_0_0_514), .B2(
      n_0_0_543), .ZN(n_0_0_548));
   OAI22_X1 i_0_0_685 (.A1(n_0_0_531), .A2(n_0_0_23), .B1(shift[2]), .B2(
      n_0_0_548), .ZN(n_0_0_549));
   AOI22_X1 i_0_0_686 (.A1(n_0_0_540), .A2(shift[1]), .B1(n_0_0_549), .B2(
      n_0_0_24), .ZN(n_0_0_550));
   OAI22_X1 i_0_0_687 (.A1(n_0_0_546), .A2(n_0_0_19), .B1(n_0_0_550), .B2(
      shift[0]), .ZN(n_0_165));
   NOR2_X1 i_0_0_688 (.A1(n_0_0_375), .A2(n_0_0_33), .ZN(n_0_0_551));
   OAI22_X1 i_0_0_689 (.A1(n_0_0_551), .A2(n_0_0_509), .B1(n_0_0_518), .B2(
      n_0_0_543), .ZN(n_0_0_552));
   OAI22_X1 i_0_0_690 (.A1(n_0_0_535), .A2(n_0_0_23), .B1(shift[2]), .B2(
      n_0_0_552), .ZN(n_0_0_553));
   AOI22_X1 i_0_0_691 (.A1(n_0_0_553), .A2(n_0_0_24), .B1(n_0_0_545), .B2(
      shift[1]), .ZN(n_0_0_554));
   OAI22_X1 i_0_0_692 (.A1(n_0_0_550), .A2(n_0_0_19), .B1(n_0_0_554), .B2(
      shift[0]), .ZN(n_0_166));
   NOR2_X1 i_0_0_693 (.A1(n_0_0_33), .A2(shift[3]), .ZN(n_0_0_555));
   AOI221_X1 i_0_0_694 (.A(n_0_0_423), .B1(n_0_0_384), .B2(n_0_0_555), .C1(
      shift[3]), .C2(n_0_0_522), .ZN(n_0_0_556));
   AOI22_X1 i_0_0_695 (.A1(n_0_0_539), .A2(shift[2]), .B1(n_0_0_556), .B2(
      n_0_0_23), .ZN(n_0_0_557));
   AOI22_X1 i_0_0_696 (.A1(n_0_0_557), .A2(n_0_0_24), .B1(n_0_0_549), .B2(
      shift[1]), .ZN(n_0_0_558));
   OAI22_X1 i_0_0_697 (.A1(n_0_0_558), .A2(shift[0]), .B1(n_0_0_554), .B2(
      n_0_0_19), .ZN(n_0_167));
   INV_X1 i_0_0_698 (.A(n_0_0_428), .ZN(n_0_0_559));
   OAI221_X1 i_0_0_699 (.A(n_0_0_295), .B1(n_0_0_392), .B2(n_0_0_428), .C1(
      n_0_0_491), .C2(n_0_0_559), .ZN(n_0_0_560));
   OAI211_X1 i_0_0_700 (.A(n_0_0_560), .B(n_0_0_23), .C1(n_0_0_526), .C2(
      n_0_0_543), .ZN(n_0_0_561));
   OAI21_X1 i_0_0_701 (.A(n_0_0_561), .B1(n_0_0_23), .B2(n_0_0_544), .ZN(
      n_0_0_562));
   AOI22_X1 i_0_0_702 (.A1(n_0_0_562), .A2(n_0_0_24), .B1(n_0_0_553), .B2(
      shift[1]), .ZN(n_0_0_563));
   OAI22_X1 i_0_0_703 (.A1(n_0_0_563), .A2(shift[0]), .B1(n_0_0_558), .B2(
      n_0_0_19), .ZN(n_0_168));
   OAI21_X1 i_0_0_704 (.A(n_0_0_23), .B1(n_0_0_530), .B2(n_0_0_543), .ZN(
      n_0_0_564));
   AOI21_X1 i_0_0_705 (.A(n_0_0_509), .B1(n_0_0_402), .B2(shift[5]), .ZN(
      n_0_0_565));
   OAI22_X1 i_0_0_706 (.A1(n_0_0_548), .A2(n_0_0_23), .B1(n_0_0_564), .B2(
      n_0_0_565), .ZN(n_0_0_566));
   OAI22_X1 i_0_0_707 (.A1(n_0_0_557), .A2(n_0_0_24), .B1(shift[1]), .B2(
      n_0_0_566), .ZN(n_0_0_567));
   OAI22_X1 i_0_0_708 (.A1(n_0_0_563), .A2(n_0_0_19), .B1(n_0_0_567), .B2(
      shift[0]), .ZN(n_0_169));
   OAI21_X1 i_0_0_709 (.A(n_0_0_23), .B1(n_0_0_534), .B2(n_0_0_543), .ZN(
      n_0_0_568));
   AOI21_X1 i_0_0_710 (.A(n_0_0_509), .B1(n_0_0_410), .B2(shift[5]), .ZN(
      n_0_0_569));
   OAI22_X1 i_0_0_711 (.A1(n_0_0_552), .A2(n_0_0_23), .B1(n_0_0_568), .B2(
      n_0_0_569), .ZN(n_0_0_570));
   OAI221_X1 i_0_0_712 (.A(n_0_0_19), .B1(shift[1]), .B2(n_0_0_570), .C1(
      n_0_0_562), .C2(n_0_0_24), .ZN(n_0_0_571));
   OAI21_X1 i_0_0_713 (.A(n_0_0_571), .B1(n_0_0_19), .B2(n_0_0_567), .ZN(n_0_170));
   DFF_X1 write_en_reg (.D(start), .CK(clk), .Q(write_en), .QN());
   DFF_X1 \c_reg[63]  (.D(n_0_104), .CK(clk), .Q(c[63]), .QN());
   DFF_X1 \c_reg[62]  (.D(n_0_103), .CK(clk), .Q(c[62]), .QN());
   DFF_X1 \c_reg[61]  (.D(n_0_102), .CK(clk), .Q(c[61]), .QN());
   DFF_X1 \c_reg[60]  (.D(n_0_101), .CK(clk), .Q(c[60]), .QN());
   DFF_X1 \c_reg[59]  (.D(n_0_100), .CK(clk), .Q(c[59]), .QN());
   DFF_X1 \c_reg[58]  (.D(n_0_99), .CK(clk), .Q(c[58]), .QN());
   DFF_X1 \c_reg[57]  (.D(n_0_98), .CK(clk), .Q(c[57]), .QN());
   DFF_X1 \c_reg[56]  (.D(n_0_97), .CK(clk), .Q(c[56]), .QN());
   DFF_X1 \c_reg[55]  (.D(n_0_96), .CK(clk), .Q(c[55]), .QN());
   DFF_X1 \c_reg[54]  (.D(n_0_95), .CK(clk), .Q(c[54]), .QN());
   DFF_X1 \c_reg[53]  (.D(n_0_94), .CK(clk), .Q(c[53]), .QN());
   DFF_X1 \c_reg[52]  (.D(n_0_93), .CK(clk), .Q(c[52]), .QN());
   DFF_X1 \c_reg[51]  (.D(n_0_92), .CK(clk), .Q(c[51]), .QN());
   DFF_X1 \c_reg[50]  (.D(n_0_91), .CK(clk), .Q(c[50]), .QN());
   DFF_X1 \c_reg[49]  (.D(n_0_90), .CK(clk), .Q(c[49]), .QN());
   DFF_X1 \c_reg[48]  (.D(n_0_89), .CK(clk), .Q(c[48]), .QN());
   DFF_X1 \c_reg[47]  (.D(n_0_88), .CK(clk), .Q(c[47]), .QN());
   DFF_X1 \c_reg[46]  (.D(n_0_87), .CK(clk), .Q(c[46]), .QN());
   DFF_X1 \c_reg[45]  (.D(n_0_86), .CK(clk), .Q(c[45]), .QN());
   DFF_X1 \c_reg[44]  (.D(n_0_85), .CK(clk), .Q(c[44]), .QN());
   DFF_X1 \c_reg[43]  (.D(n_0_84), .CK(clk), .Q(c[43]), .QN());
   DFF_X1 \c_reg[42]  (.D(n_0_83), .CK(clk), .Q(c[42]), .QN());
   DFF_X1 \c_reg[41]  (.D(n_0_82), .CK(clk), .Q(c[41]), .QN());
   DFF_X1 \c_reg[40]  (.D(n_0_81), .CK(clk), .Q(c[40]), .QN());
   DFF_X1 \c_reg[39]  (.D(n_0_80), .CK(clk), .Q(c[39]), .QN());
   DFF_X1 \c_reg[38]  (.D(n_0_79), .CK(clk), .Q(c[38]), .QN());
   DFF_X1 \c_reg[37]  (.D(n_0_78), .CK(clk), .Q(c[37]), .QN());
   DFF_X1 \c_reg[36]  (.D(n_0_77), .CK(clk), .Q(c[36]), .QN());
   DFF_X1 \c_reg[35]  (.D(n_0_76), .CK(clk), .Q(c[35]), .QN());
   DFF_X1 \c_reg[34]  (.D(n_0_269), .CK(clk), .Q(c[34]), .QN());
   DFF_X1 \c_reg[33]  (.D(n_0_268), .CK(clk), .Q(c[33]), .QN());
   DFF_X1 \c_reg[32]  (.D(n_0_267), .CK(clk), .Q(c[32]), .QN());
   DFF_X1 \c_reg[31]  (.D(n_0_266), .CK(clk), .Q(c[31]), .QN());
   DFF_X1 \c_reg[30]  (.D(n_0_265), .CK(clk), .Q(c[30]), .QN());
   DFF_X1 \c_reg[29]  (.D(n_0_264), .CK(clk), .Q(c[29]), .QN());
   DFF_X1 \c_reg[28]  (.D(n_0_263), .CK(clk), .Q(c[28]), .QN());
   DFF_X1 \c_reg[27]  (.D(n_0_262), .CK(clk), .Q(c[27]), .QN());
   DFF_X1 \c_reg[26]  (.D(n_0_261), .CK(clk), .Q(c[26]), .QN());
   DFF_X1 \c_reg[25]  (.D(n_0_260), .CK(clk), .Q(c[25]), .QN());
   DFF_X1 \c_reg[24]  (.D(n_0_259), .CK(clk), .Q(c[24]), .QN());
   DFF_X1 \c_reg[23]  (.D(n_0_258), .CK(clk), .Q(c[23]), .QN());
   DFF_X1 \c_reg[22]  (.D(n_0_257), .CK(clk), .Q(c[22]), .QN());
   DFF_X1 \c_reg[21]  (.D(n_0_256), .CK(clk), .Q(c[21]), .QN());
   DFF_X1 \c_reg[20]  (.D(n_0_255), .CK(clk), .Q(c[20]), .QN());
   DFF_X1 \c_reg[19]  (.D(n_0_254), .CK(clk), .Q(c[19]), .QN());
   DFF_X1 \c_reg[18]  (.D(n_0_253), .CK(clk), .Q(c[18]), .QN());
   DFF_X1 \c_reg[17]  (.D(n_0_252), .CK(clk), .Q(c[17]), .QN());
   DFF_X1 \c_reg[16]  (.D(n_0_251), .CK(clk), .Q(c[16]), .QN());
   DFF_X1 \c_reg[15]  (.D(n_0_250), .CK(clk), .Q(c[15]), .QN());
   DFF_X1 \c_reg[14]  (.D(n_0_249), .CK(clk), .Q(c[14]), .QN());
   DFF_X1 \c_reg[13]  (.D(n_0_248), .CK(clk), .Q(c[13]), .QN());
   DFF_X1 \c_reg[12]  (.D(n_0_247), .CK(clk), .Q(c[12]), .QN());
   DFF_X1 \c_reg[11]  (.D(n_0_246), .CK(clk), .Q(c[11]), .QN());
   DFF_X1 \c_reg[10]  (.D(n_0_245), .CK(clk), .Q(c[10]), .QN());
   DFF_X1 \c_reg[9]  (.D(n_0_244), .CK(clk), .Q(c[9]), .QN());
   DFF_X1 \c_reg[8]  (.D(n_0_243), .CK(clk), .Q(c[8]), .QN());
   DFF_X1 \c_reg[7]  (.D(n_0_242), .CK(clk), .Q(c[7]), .QN());
   DFF_X1 \c_reg[6]  (.D(n_0_241), .CK(clk), .Q(c[6]), .QN());
   DFF_X1 \c_reg[5]  (.D(n_0_240), .CK(clk), .Q(c[5]), .QN());
   DFF_X1 \c_reg[4]  (.D(n_0_239), .CK(clk), .Q(c[4]), .QN());
   DFF_X1 \c_reg[3]  (.D(n_0_238), .CK(clk), .Q(c[3]), .QN());
   DFF_X1 \c_reg[2]  (.D(n_0_237), .CK(clk), .Q(c[2]), .QN());
   DFF_X1 \c_reg[1]  (.D(n_0_236), .CK(clk), .Q(c[1]), .QN());
   DFF_X1 \c_reg[0]  (.D(n_0_235), .CK(clk), .Q(c[0]), .QN());
   DFF_X1 \shift_reg[5]  (.D(n_0_75), .CK(n_0_106), .Q(shift[5]), .QN());
   DFF_X1 \shift_reg[4]  (.D(n_0_74), .CK(n_0_106), .Q(shift[4]), .QN());
   DFF_X1 \shift_reg[3]  (.D(n_0_73), .CK(n_0_106), .Q(shift[3]), .QN());
   DFF_X1 \shift_reg[2]  (.D(n_0_72), .CK(n_0_106), .Q(shift[2]), .QN());
   DFF_X1 \shift_reg[1]  (.D(n_0_71), .CK(n_0_106), .Q(shift[1]), .QN());
   DFF_X1 \shift_reg[0]  (.D(n_0_70), .CK(n_0_106), .Q(shift[0]), .QN());
   DFF_X1 \i_reg[5]  (.D(n_0_68), .CK(n_0_106), .Q(i[5]), .QN());
   DFF_X1 \i_reg[4]  (.D(n_0_67), .CK(n_0_106), .Q(i[4]), .QN());
   DFF_X1 \i_reg[3]  (.D(n_0_66), .CK(n_0_106), .Q(i[3]), .QN());
   DFF_X1 \i_reg[2]  (.D(n_0_3), .CK(n_0_106), .Q(i[2]), .QN());
   DFF_X1 \i_reg[1]  (.D(n_0_2), .CK(n_0_106), .Q(i[1]), .QN());
   DFF_X1 \i_reg[0]  (.D(n_0_1), .CK(n_0_106), .Q(i[0]), .QN());
   CLKGATETST_X1 clk_gate_i_reg (.CK(clk), .E(n_0_69), .SE(1'b0), .GCK(n_0_106));
endmodule
