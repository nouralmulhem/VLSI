
// 	Sat Dec 24 09:10:58 2022
//	vlsi
//	localhost.localdomain

module datapath__0_17 (f8, p_0);

output [31:0] p_0;
input [31:0] f8;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (f8[25]));
INV_X1 i_63 (.ZN (n_32), .A (f8[21]));
INV_X1 i_62 (.ZN (n_31), .A (f8[14]));
INV_X1 i_61 (.ZN (n_30), .A (f8[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (f8[2]), .A2 (f8[1]), .A3 (f8[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (f8[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (f8[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (f8[5]), .A3 (f8[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (f8[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (f8[8]), .A3 (f8[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (f8[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (f8[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (f8[12]), .A3 (f8[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (f8[15]), .A3 (f8[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (f8[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (f8[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (f8[18]), .A3 (f8[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (f8[18]), .A3 (f8[19]), .A4 (f8[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (f8[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (f8[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (f8[23]), .A3 (f8[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (f8[26]), .A3 (f8[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (f8[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (f8[28]), .A3 (f8[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (f8[28]), .A3 (f8[29]), .A4 (f8[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (f8[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (f8[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (f8[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (f8[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (f8[27]), .B1 (n_9), .B2 (f8[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (f8[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (f8[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (f8[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (f8[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (f8[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (f8[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (f8[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (f8[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (f8[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (f8[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (f8[16]), .B1 (n_19), .B2 (f8[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (f8[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (f8[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (f8[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (f8[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (f8[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (f8[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (f8[9]), .B1 (n_25), .B2 (f8[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (f8[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (f8[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (f8[6]), .B1 (n_27), .B2 (f8[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (f8[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (f8[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (f8[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (f8[2]), .B1 (f8[1]), .B2 (f8[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (f8[1]), .B (f8[0]));

endmodule //datapath__0_17

module regFile (clk_CTS_1_PP_0, read_data, read_data2, write_en, write_data, write_data2, 
    clk);

output [31:0] read_data2;
output [31:0] read_data;
input clk;
input [31:0] write_data2;
input [31:0] write_data;
input write_en;
input clk_CTS_1_PP_0;
wire CTS_n_tid1_2;
wire CTS_n_tid1_3;


CLKGATETST_X8 clk_gate_my_reg_reg (.GCK (CTS_n_tid1_3), .CK (clk_CTS_1_PP_0), .E (write_en), .SE (1'b0 ));
DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid1_2), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid1_2), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid1_2), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid1_2), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid1_2), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid1_2), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid1_2), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid1_2), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid1_2), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid1_2), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid1_2), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid1_2), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid1_2), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid1_2), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid1_2), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid1_2), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid1_2), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid1_2), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid1_2), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid1_2), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid1_2), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid1_2), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid1_2), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid1_2), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid1_2), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid1_2), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid1_2), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid1_2), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid1_2), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid1_2), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid1_2), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid1_2), .D (write_data[31]));
DFF_X1 \my_reg2_reg[0]  (.Q (read_data2[0]), .CK (CTS_n_tid1_2), .D (write_data2[0]));
DFF_X1 \my_reg2_reg[1]  (.Q (read_data2[1]), .CK (CTS_n_tid1_2), .D (write_data2[1]));
DFF_X1 \my_reg2_reg[2]  (.Q (read_data2[2]), .CK (CTS_n_tid1_2), .D (write_data2[2]));
DFF_X1 \my_reg2_reg[3]  (.Q (read_data2[3]), .CK (CTS_n_tid1_2), .D (write_data2[3]));
DFF_X1 \my_reg2_reg[4]  (.Q (read_data2[4]), .CK (CTS_n_tid1_2), .D (write_data2[4]));
DFF_X1 \my_reg2_reg[5]  (.Q (read_data2[5]), .CK (CTS_n_tid1_2), .D (write_data2[5]));
DFF_X1 \my_reg2_reg[6]  (.Q (read_data2[6]), .CK (CTS_n_tid1_2), .D (write_data2[6]));
DFF_X1 \my_reg2_reg[7]  (.Q (read_data2[7]), .CK (CTS_n_tid1_2), .D (write_data2[7]));
DFF_X1 \my_reg2_reg[8]  (.Q (read_data2[8]), .CK (CTS_n_tid1_2), .D (write_data2[8]));
DFF_X1 \my_reg2_reg[9]  (.Q (read_data2[9]), .CK (CTS_n_tid1_2), .D (write_data2[9]));
DFF_X1 \my_reg2_reg[10]  (.Q (read_data2[10]), .CK (CTS_n_tid1_2), .D (write_data2[10]));
DFF_X1 \my_reg2_reg[11]  (.Q (read_data2[11]), .CK (CTS_n_tid1_2), .D (write_data2[11]));
DFF_X1 \my_reg2_reg[12]  (.Q (read_data2[12]), .CK (CTS_n_tid1_2), .D (write_data2[12]));
DFF_X1 \my_reg2_reg[13]  (.Q (read_data2[13]), .CK (CTS_n_tid1_2), .D (write_data2[13]));
DFF_X1 \my_reg2_reg[14]  (.Q (read_data2[14]), .CK (CTS_n_tid1_2), .D (write_data2[14]));
DFF_X1 \my_reg2_reg[15]  (.Q (read_data2[15]), .CK (CTS_n_tid1_2), .D (write_data2[15]));
DFF_X1 \my_reg2_reg[16]  (.Q (read_data2[16]), .CK (CTS_n_tid1_2), .D (write_data2[16]));
DFF_X1 \my_reg2_reg[17]  (.Q (read_data2[17]), .CK (CTS_n_tid1_2), .D (write_data2[17]));
DFF_X1 \my_reg2_reg[18]  (.Q (read_data2[18]), .CK (CTS_n_tid1_2), .D (write_data2[18]));
DFF_X1 \my_reg2_reg[19]  (.Q (read_data2[19]), .CK (CTS_n_tid1_2), .D (write_data2[19]));
DFF_X1 \my_reg2_reg[20]  (.Q (read_data2[20]), .CK (CTS_n_tid1_2), .D (write_data2[20]));
DFF_X1 \my_reg2_reg[21]  (.Q (read_data2[21]), .CK (CTS_n_tid1_2), .D (write_data2[21]));
DFF_X1 \my_reg2_reg[22]  (.Q (read_data2[22]), .CK (CTS_n_tid1_2), .D (write_data2[22]));
DFF_X1 \my_reg2_reg[23]  (.Q (read_data2[23]), .CK (CTS_n_tid1_2), .D (write_data2[23]));
DFF_X1 \my_reg2_reg[24]  (.Q (read_data2[24]), .CK (CTS_n_tid1_2), .D (write_data2[24]));
DFF_X1 \my_reg2_reg[25]  (.Q (read_data2[25]), .CK (CTS_n_tid1_2), .D (write_data2[25]));
DFF_X1 \my_reg2_reg[26]  (.Q (read_data2[26]), .CK (CTS_n_tid1_2), .D (write_data2[26]));
DFF_X1 \my_reg2_reg[27]  (.Q (read_data2[27]), .CK (CTS_n_tid1_2), .D (write_data2[27]));
DFF_X1 \my_reg2_reg[28]  (.Q (read_data2[28]), .CK (CTS_n_tid1_2), .D (write_data2[28]));
DFF_X1 \my_reg2_reg[29]  (.Q (read_data2[29]), .CK (CTS_n_tid1_2), .D (write_data2[29]));
DFF_X1 \my_reg2_reg[30]  (.Q (read_data2[30]), .CK (CTS_n_tid1_2), .D (write_data2[30]));
DFF_X1 \my_reg2_reg[31]  (.Q (read_data2[31]), .CK (CTS_n_tid1_2), .D (write_data2[31]));
CLKBUF_X3 CTS_L3_c_tid1_3 (.Z (CTS_n_tid1_2), .A (CTS_n_tid1_3));

endmodule //regFile

module fullAdder (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (y));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (x), .B (cin));

endmodule //fullAdder

module fullAdder__0_207 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_207

module fullAdder__0_204 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_204

module fullAdder__0_201 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_201

module fullAdder__0_198 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_198

module fullAdder__0_195 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_195

module fullAdder__0_192 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_192

module fullAdder__0_189 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_189

module fullAdder__0_186 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_186

module fullAdder__0_183 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_183

module fullAdder__0_180 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_180

module fullAdder__0_177 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_177

module fullAdder__0_174 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_174

module fullAdder__0_171 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_171

module fullAdder__0_168 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_168

module fullAdder__0_165 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_165

module fullAdder__0_162 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_162

module fullAdder__0_159 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_159

module fullAdder__0_156 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_156

module fullAdder__0_153 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_153

module fullAdder__0_150 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_150

module fullAdder__0_147 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_147

module fullAdder__0_144 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_144

module fullAdder__0_141 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_141

module fullAdder__0_138 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_138

module fullAdder__0_135 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_135

module fullAdder__0_132 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_132

module fullAdder__0_129 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_129

module fullAdder__0_126 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_126

module fullAdder__0_123 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_123

module fullAdder__0_120 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


XOR2_X1 i_0_0 (.Z (sum), .A (y), .B (x));

endmodule //fullAdder__0_120

module fullAdder__0_117 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_117

module fullAdder__0_114 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_114

module fullAdder__0_111 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_111

module fullAdder__0_108 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_108

module fullAdder__0_105 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_105

module fullAdder__0_102 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_102

module fullAdder__0_99 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_99

module fullAdder__0_96 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_96

module fullAdder__0_93 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_93

module fullAdder__0_90 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_90

module fullAdder__0_87 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_87

module fullAdder__0_84 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_84

module fullAdder__0_81 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_81

module fullAdder__0_78 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_78

module fullAdder__0_75 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_75

module fullAdder__0_72 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_72

module fullAdder__0_69 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_69

module fullAdder__0_66 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_66

module fullAdder__0_63 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_63

module fullAdder__0_60 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_60

module fullAdder__0_57 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_57

module fullAdder__0_54 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_54

module fullAdder__0_51 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_51

module fullAdder__0_48 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_48

module fullAdder__0_45 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_45

module fullAdder__0_42 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_42

module fullAdder__0_39 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_39

module fullAdder__0_36 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_36

module fullAdder__0_33 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_33

module fullAdder__0_30 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_30

module fullAdder__0_27 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_27

module fullAdder__0_21 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_21

module carrySaveAdder (a, b, c, sum, cout);

output cout;
output [31:0] sum;
input [31:0] a;
input [31:0] b;
input [31:0] c;
wire \halfcarry[29] ;
wire \halfcarry[28] ;
wire \halfcarry[27] ;
wire \halfcarry[26] ;
wire \halfcarry[25] ;
wire \halfcarry[24] ;
wire \halfcarry[23] ;
wire \halfcarry[22] ;
wire \halfcarry[21] ;
wire \halfcarry[20] ;
wire \halfcarry[19] ;
wire \halfcarry[18] ;
wire \halfcarry[17] ;
wire \halfcarry[16] ;
wire \halfcarry[15] ;
wire \halfcarry[14] ;
wire \halfcarry[13] ;
wire \halfcarry[12] ;
wire \halfcarry[11] ;
wire \halfcarry[10] ;
wire \halfcarry[9] ;
wire \halfcarry[8] ;
wire \halfcarry[7] ;
wire \halfcarry[6] ;
wire \halfcarry[5] ;
wire \halfcarry[4] ;
wire \halfcarry[3] ;
wire \halfcarry[2] ;
wire \halfcarry[1] ;
wire \halfcarry[0] ;
wire \halfcout[30] ;
wire \halfcout[29] ;
wire \halfcout[28] ;
wire \halfcout[27] ;
wire \halfcout[26] ;
wire \halfcout[25] ;
wire \halfcout[24] ;
wire \halfcout[23] ;
wire \halfcout[22] ;
wire \halfcout[21] ;
wire \halfcout[20] ;
wire \halfcout[19] ;
wire \halfcout[18] ;
wire \halfcout[17] ;
wire \halfcout[16] ;
wire \halfcout[15] ;
wire \halfcout[14] ;
wire \halfcout[13] ;
wire \halfcout[12] ;
wire \halfcout[11] ;
wire \halfcout[10] ;
wire \halfcout[9] ;
wire \halfcout[8] ;
wire \halfcout[7] ;
wire \halfcout[6] ;
wire \halfcout[5] ;
wire \halfcout[4] ;
wire \halfcout[3] ;
wire \halfcout[2] ;
wire \halfcout[1] ;
wire \halfcout[0] ;
wire \halfsum[31] ;
wire \halfsum[30] ;
wire \halfsum[29] ;
wire \halfsum[28] ;
wire \halfsum[27] ;
wire \halfsum[26] ;
wire \halfsum[25] ;
wire \halfsum[24] ;
wire \halfsum[23] ;
wire \halfsum[22] ;
wire \halfsum[21] ;
wire \halfsum[20] ;
wire \halfsum[19] ;
wire \halfsum[18] ;
wire \halfsum[17] ;
wire \halfsum[16] ;
wire \halfsum[15] ;
wire \halfsum[14] ;
wire \halfsum[13] ;
wire \halfsum[12] ;
wire \halfsum[11] ;
wire \halfsum[10] ;
wire \halfsum[9] ;
wire \halfsum[8] ;
wire \halfsum[7] ;
wire \halfsum[6] ;
wire \halfsum[5] ;
wire \halfsum[4] ;
wire \halfsum[3] ;
wire \halfsum[2] ;
wire \halfsum[1] ;


fullAdder genblk2_30_f3 (.sum (sum[31]), .cin (\halfcarry[29] ), .x (\halfsum[31] ), .y (\halfcout[30] ));
fullAdder__0_207 genblk2_29_f3 (.cout (\halfcarry[29] ), .sum (sum[30]), .cin (\halfcarry[28] )
    , .x (\halfsum[30] ), .y (\halfcout[29] ));
fullAdder__0_204 genblk2_28_f3 (.cout (\halfcarry[28] ), .sum (sum[29]), .cin (\halfcarry[27] )
    , .x (\halfsum[29] ), .y (\halfcout[28] ));
fullAdder__0_201 genblk2_27_f3 (.cout (\halfcarry[27] ), .sum (sum[28]), .cin (\halfcarry[26] )
    , .x (\halfsum[28] ), .y (\halfcout[27] ));
fullAdder__0_198 genblk2_26_f3 (.cout (\halfcarry[26] ), .sum (sum[27]), .cin (\halfcarry[25] )
    , .x (\halfsum[27] ), .y (\halfcout[26] ));
fullAdder__0_195 genblk2_25_f3 (.cout (\halfcarry[25] ), .sum (sum[26]), .cin (\halfcarry[24] )
    , .x (\halfsum[26] ), .y (\halfcout[25] ));
fullAdder__0_192 genblk2_24_f3 (.cout (\halfcarry[24] ), .sum (sum[25]), .cin (\halfcarry[23] )
    , .x (\halfsum[25] ), .y (\halfcout[24] ));
fullAdder__0_189 genblk2_23_f3 (.cout (\halfcarry[23] ), .sum (sum[24]), .cin (\halfcarry[22] )
    , .x (\halfsum[24] ), .y (\halfcout[23] ));
fullAdder__0_186 genblk2_22_f3 (.cout (\halfcarry[22] ), .sum (sum[23]), .cin (\halfcarry[21] )
    , .x (\halfsum[23] ), .y (\halfcout[22] ));
fullAdder__0_183 genblk2_21_f3 (.cout (\halfcarry[21] ), .sum (sum[22]), .cin (\halfcarry[20] )
    , .x (\halfsum[22] ), .y (\halfcout[21] ));
fullAdder__0_180 genblk2_20_f3 (.cout (\halfcarry[20] ), .sum (sum[21]), .cin (\halfcarry[19] )
    , .x (\halfsum[21] ), .y (\halfcout[20] ));
fullAdder__0_177 genblk2_19_f3 (.cout (\halfcarry[19] ), .sum (sum[20]), .cin (\halfcarry[18] )
    , .x (\halfsum[20] ), .y (\halfcout[19] ));
fullAdder__0_174 genblk2_18_f3 (.cout (\halfcarry[18] ), .sum (sum[19]), .cin (\halfcarry[17] )
    , .x (\halfsum[19] ), .y (\halfcout[18] ));
fullAdder__0_171 genblk2_17_f3 (.cout (\halfcarry[17] ), .sum (sum[18]), .cin (\halfcarry[16] )
    , .x (\halfsum[18] ), .y (\halfcout[17] ));
fullAdder__0_168 genblk2_16_f3 (.cout (\halfcarry[16] ), .sum (sum[17]), .cin (\halfcarry[15] )
    , .x (\halfsum[17] ), .y (\halfcout[16] ));
fullAdder__0_165 genblk2_15_f3 (.cout (\halfcarry[15] ), .sum (sum[16]), .cin (\halfcarry[14] )
    , .x (\halfsum[16] ), .y (\halfcout[15] ));
fullAdder__0_162 genblk2_14_f3 (.cout (\halfcarry[14] ), .sum (sum[15]), .cin (\halfcarry[13] )
    , .x (\halfsum[15] ), .y (\halfcout[14] ));
fullAdder__0_159 genblk2_13_f3 (.cout (\halfcarry[13] ), .sum (sum[14]), .cin (\halfcarry[12] )
    , .x (\halfsum[14] ), .y (\halfcout[13] ));
fullAdder__0_156 genblk2_12_f3 (.cout (\halfcarry[12] ), .sum (sum[13]), .cin (\halfcarry[11] )
    , .x (\halfsum[13] ), .y (\halfcout[12] ));
fullAdder__0_153 genblk2_11_f3 (.cout (\halfcarry[11] ), .sum (sum[12]), .cin (\halfcarry[10] )
    , .x (\halfsum[12] ), .y (\halfcout[11] ));
fullAdder__0_150 genblk2_10_f3 (.cout (\halfcarry[10] ), .sum (sum[11]), .cin (\halfcarry[9] )
    , .x (\halfsum[11] ), .y (\halfcout[10] ));
fullAdder__0_147 genblk2_9_f3 (.cout (\halfcarry[9] ), .sum (sum[10]), .cin (\halfcarry[8] )
    , .x (\halfsum[10] ), .y (\halfcout[9] ));
fullAdder__0_144 genblk2_8_f3 (.cout (\halfcarry[8] ), .sum (sum[9]), .cin (\halfcarry[7] )
    , .x (\halfsum[9] ), .y (\halfcout[8] ));
fullAdder__0_141 genblk2_7_f3 (.cout (\halfcarry[7] ), .sum (sum[8]), .cin (\halfcarry[6] )
    , .x (\halfsum[8] ), .y (\halfcout[7] ));
fullAdder__0_138 genblk2_6_f3 (.cout (\halfcarry[6] ), .sum (sum[7]), .cin (\halfcarry[5] )
    , .x (\halfsum[7] ), .y (\halfcout[6] ));
fullAdder__0_135 genblk2_5_f3 (.cout (\halfcarry[5] ), .sum (sum[6]), .cin (\halfcarry[4] )
    , .x (\halfsum[6] ), .y (\halfcout[5] ));
fullAdder__0_132 genblk2_4_f3 (.cout (\halfcarry[4] ), .sum (sum[5]), .cin (\halfcarry[3] )
    , .x (\halfsum[5] ), .y (\halfcout[4] ));
fullAdder__0_129 genblk2_3_f3 (.cout (\halfcarry[3] ), .sum (sum[4]), .cin (\halfcarry[2] )
    , .x (\halfsum[4] ), .y (\halfcout[3] ));
fullAdder__0_126 genblk2_2_f3 (.cout (\halfcarry[2] ), .sum (sum[3]), .cin (\halfcarry[1] )
    , .x (\halfsum[3] ), .y (\halfcout[2] ));
fullAdder__0_123 genblk2_1_f3 (.cout (\halfcarry[1] ), .sum (sum[2]), .cin (\halfcarry[0] )
    , .x (\halfsum[2] ), .y (\halfcout[1] ));
fullAdder__0_120 genblk1_31_fulladder_f1 (.sum (\halfsum[31] ), .x (a[31]), .y (b[31]));
fullAdder__0_117 genblk1_30_fulladder_f1 (.cout (\halfcout[30] ), .sum (\halfsum[30] )
    , .x (a[30]), .y (b[30]));
fullAdder__0_114 genblk1_29_fulladder_f1 (.cout (\halfcout[29] ), .sum (\halfsum[29] )
    , .x (a[29]), .y (b[29]));
fullAdder__0_111 genblk1_28_fulladder_f1 (.cout (\halfcout[28] ), .sum (\halfsum[28] )
    , .x (a[28]), .y (b[28]));
fullAdder__0_108 genblk1_27_fulladder_f1 (.cout (\halfcout[27] ), .sum (\halfsum[27] )
    , .x (a[27]), .y (b[27]));
fullAdder__0_105 genblk1_26_fulladder_f1 (.cout (\halfcout[26] ), .sum (\halfsum[26] )
    , .x (a[26]), .y (b[26]));
fullAdder__0_102 genblk1_25_fulladder_f1 (.cout (\halfcout[25] ), .sum (\halfsum[25] )
    , .x (a[25]), .y (b[25]));
fullAdder__0_99 genblk1_24_fulladder_f1 (.cout (\halfcout[24] ), .sum (\halfsum[24] )
    , .x (a[24]), .y (b[24]));
fullAdder__0_96 genblk1_23_fulladder_f1 (.cout (\halfcout[23] ), .sum (\halfsum[23] )
    , .x (a[23]), .y (b[23]));
fullAdder__0_93 genblk1_22_fulladder_f1 (.cout (\halfcout[22] ), .sum (\halfsum[22] )
    , .x (a[22]), .y (b[22]));
fullAdder__0_90 genblk1_21_fulladder_f1 (.cout (\halfcout[21] ), .sum (\halfsum[21] )
    , .x (a[21]), .y (b[21]));
fullAdder__0_87 genblk1_20_fulladder_f1 (.cout (\halfcout[20] ), .sum (\halfsum[20] )
    , .x (a[20]), .y (b[20]));
fullAdder__0_84 genblk1_19_fulladder_f1 (.cout (\halfcout[19] ), .sum (\halfsum[19] )
    , .x (a[19]), .y (b[19]));
fullAdder__0_81 genblk1_18_fulladder_f1 (.cout (\halfcout[18] ), .sum (\halfsum[18] )
    , .x (a[18]), .y (b[18]));
fullAdder__0_78 genblk1_17_fulladder_f1 (.cout (\halfcout[17] ), .sum (\halfsum[17] )
    , .x (a[17]), .y (b[17]));
fullAdder__0_75 genblk1_16_fulladder_f1 (.cout (\halfcout[16] ), .sum (\halfsum[16] )
    , .x (a[16]), .y (b[16]));
fullAdder__0_72 genblk1_15_fulladder_f1 (.cout (\halfcout[15] ), .sum (\halfsum[15] )
    , .x (a[15]), .y (b[15]));
fullAdder__0_69 genblk1_14_fulladder_f1 (.cout (\halfcout[14] ), .sum (\halfsum[14] )
    , .x (a[14]), .y (b[14]));
fullAdder__0_66 genblk1_13_fulladder_f1 (.cout (\halfcout[13] ), .sum (\halfsum[13] )
    , .x (a[13]), .y (b[13]));
fullAdder__0_63 genblk1_12_fulladder_f1 (.cout (\halfcout[12] ), .sum (\halfsum[12] )
    , .x (a[12]), .y (b[12]));
fullAdder__0_60 genblk1_11_fulladder_f1 (.cout (\halfcout[11] ), .sum (\halfsum[11] )
    , .x (a[11]), .y (b[11]));
fullAdder__0_57 genblk1_10_fulladder_f1 (.cout (\halfcout[10] ), .sum (\halfsum[10] )
    , .x (a[10]), .y (b[10]));
fullAdder__0_54 genblk1_9_fulladder_f1 (.cout (\halfcout[9] ), .sum (\halfsum[9] )
    , .x (a[9]), .y (b[9]));
fullAdder__0_51 genblk1_8_fulladder_f1 (.cout (\halfcout[8] ), .sum (\halfsum[8] )
    , .x (a[8]), .y (b[8]));
fullAdder__0_48 genblk1_7_fulladder_f1 (.cout (\halfcout[7] ), .sum (\halfsum[7] )
    , .x (a[7]), .y (b[7]));
fullAdder__0_45 genblk1_6_fulladder_f1 (.cout (\halfcout[6] ), .sum (\halfsum[6] )
    , .x (a[6]), .y (b[6]));
fullAdder__0_42 genblk1_5_fulladder_f1 (.cout (\halfcout[5] ), .sum (\halfsum[5] )
    , .x (a[5]), .y (b[5]));
fullAdder__0_39 genblk1_4_fulladder_f1 (.cout (\halfcout[4] ), .sum (\halfsum[4] )
    , .x (a[4]), .y (b[4]));
fullAdder__0_36 genblk1_3_fulladder_f1 (.cout (\halfcout[3] ), .sum (\halfsum[3] )
    , .x (a[3]), .y (b[3]));
fullAdder__0_33 genblk1_2_fulladder_f1 (.cout (\halfcout[2] ), .sum (\halfsum[2] )
    , .x (a[2]), .y (b[2]));
fullAdder__0_30 genblk1_1_fulladder_f1 (.cout (\halfcout[1] ), .sum (\halfsum[1] )
    , .x (a[1]), .y (b[1]));
fullAdder__0_27 genblk1_0_fulladder_f1 (.cout (\halfcout[0] ), .sum (sum[0]), .x (a[0]), .y (b[0]));
fullAdder__0_21 fulladder_f2 (.cout (\halfcarry[0] ), .sum (sum[1]), .x (\halfsum[1] ), .y (\halfcout[0] ));

endmodule //carrySaveAdder

module fullAdder__0_210 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;


XNOR2_X1 i_0_1 (.ZN (sum), .A (n_0_0), .B (y));
XNOR2_X1 i_0_0 (.ZN (n_0_0), .A (x), .B (cin));

endmodule //fullAdder__0_210

module fullAdder__0_213 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_213

module fullAdder__0_216 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_216

module fullAdder__0_219 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_219

module fullAdder__0_222 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_222

module fullAdder__0_225 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_225

module fullAdder__0_228 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_228

module fullAdder__0_231 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_231

module fullAdder__0_234 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_234

module fullAdder__0_237 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_237

module fullAdder__0_240 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_240

module fullAdder__0_243 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_243

module fullAdder__0_246 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_246

module fullAdder__0_249 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_249

module fullAdder__0_252 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_252

module fullAdder__0_255 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_255

module fullAdder__0_258 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_258

module fullAdder__0_261 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_261

module fullAdder__0_264 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_264

module fullAdder__0_267 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_267

module fullAdder__0_270 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_270

module fullAdder__0_273 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_273

module fullAdder__0_276 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_276

module fullAdder__0_279 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_279

module fullAdder__0_282 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_282

module fullAdder__0_285 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_285

module fullAdder__0_288 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_288

module fullAdder__0_291 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_291

module fullAdder__0_294 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_294

module fullAdder__0_297 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (cin), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (cin), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (y), .B1 (cin), .B2 (x));
NAND2_X1 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //fullAdder__0_297

module fullAdder__0_300 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


XOR2_X1 i_0_0 (.Z (sum), .A (y), .B (x));

endmodule //fullAdder__0_300

module fullAdder__0_303 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_303

module fullAdder__0_306 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_306

module fullAdder__0_309 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_309

module fullAdder__0_312 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_312

module fullAdder__0_315 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_315

module fullAdder__0_318 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_318

module fullAdder__0_321 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_321

module fullAdder__0_324 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_324

module fullAdder__0_327 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_327

module fullAdder__0_330 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_330

module fullAdder__0_333 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_333

module fullAdder__0_336 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_336

module fullAdder__0_339 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_339

module fullAdder__0_342 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_342

module fullAdder__0_345 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_345

module fullAdder__0_348 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_348

module fullAdder__0_351 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_351

module fullAdder__0_354 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_354

module fullAdder__0_357 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_357

module fullAdder__0_360 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_360

module fullAdder__0_363 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_363

module fullAdder__0_366 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_366

module fullAdder__0_369 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_369

module fullAdder__0_372 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_372

module fullAdder__0_375 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_375

module fullAdder__0_378 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_378

module fullAdder__0_381 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_381

module fullAdder__0_384 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_384

module fullAdder__0_387 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_387

module fullAdder__0_390 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_390

module fullAdder__0_393 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_393

module fullAdder__0_399 (x, y, cin, sum, cout);

output cout;
output sum;
input cin;
input x;
input y;


AND2_X1 i_0_1 (.ZN (cout), .A1 (y), .A2 (x));
XOR2_X1 i_0_0 (.Z (sum), .A (x), .B (y));

endmodule //fullAdder__0_399

module carrySaveAdder__0_400 (a, b, c, sum, cout);

output cout;
output [31:0] sum;
input [31:0] a;
input [31:0] b;
input [31:0] c;
wire \halfcarry[29] ;
wire \halfcarry[28] ;
wire \halfcarry[27] ;
wire \halfcarry[26] ;
wire \halfcarry[25] ;
wire \halfcarry[24] ;
wire \halfcarry[23] ;
wire \halfcarry[22] ;
wire \halfcarry[21] ;
wire \halfcarry[20] ;
wire \halfcarry[19] ;
wire \halfcarry[18] ;
wire \halfcarry[17] ;
wire \halfcarry[16] ;
wire \halfcarry[15] ;
wire \halfcarry[14] ;
wire \halfcarry[13] ;
wire \halfcarry[12] ;
wire \halfcarry[11] ;
wire \halfcarry[10] ;
wire \halfcarry[9] ;
wire \halfcarry[8] ;
wire \halfcarry[7] ;
wire \halfcarry[6] ;
wire \halfcarry[5] ;
wire \halfcarry[4] ;
wire \halfcarry[3] ;
wire \halfcarry[2] ;
wire \halfcarry[1] ;
wire \halfcarry[0] ;
wire \halfcout[30] ;
wire \halfcout[29] ;
wire \halfcout[28] ;
wire \halfcout[27] ;
wire \halfcout[26] ;
wire \halfcout[25] ;
wire \halfcout[24] ;
wire \halfcout[23] ;
wire \halfcout[22] ;
wire \halfcout[21] ;
wire \halfcout[20] ;
wire \halfcout[19] ;
wire \halfcout[18] ;
wire \halfcout[17] ;
wire \halfcout[16] ;
wire \halfcout[15] ;
wire \halfcout[14] ;
wire \halfcout[13] ;
wire \halfcout[12] ;
wire \halfcout[11] ;
wire \halfcout[10] ;
wire \halfcout[9] ;
wire \halfcout[8] ;
wire \halfcout[7] ;
wire \halfcout[6] ;
wire \halfcout[5] ;
wire \halfcout[4] ;
wire \halfcout[3] ;
wire \halfcout[2] ;
wire \halfcout[1] ;
wire \halfcout[0] ;
wire \halfsum[31] ;
wire \halfsum[30] ;
wire \halfsum[29] ;
wire \halfsum[28] ;
wire \halfsum[27] ;
wire \halfsum[26] ;
wire \halfsum[25] ;
wire \halfsum[24] ;
wire \halfsum[23] ;
wire \halfsum[22] ;
wire \halfsum[21] ;
wire \halfsum[20] ;
wire \halfsum[19] ;
wire \halfsum[18] ;
wire \halfsum[17] ;
wire \halfsum[16] ;
wire \halfsum[15] ;
wire \halfsum[14] ;
wire \halfsum[13] ;
wire \halfsum[12] ;
wire \halfsum[11] ;
wire \halfsum[10] ;
wire \halfsum[9] ;
wire \halfsum[8] ;
wire \halfsum[7] ;
wire \halfsum[6] ;
wire \halfsum[5] ;
wire \halfsum[4] ;
wire \halfsum[3] ;
wire \halfsum[2] ;
wire \halfsum[1] ;


fullAdder__0_210 genblk2_30_f3 (.sum (sum[31]), .cin (\halfcarry[29] ), .x (\halfsum[31] ), .y (\halfcout[30] ));
fullAdder__0_213 genblk2_29_f3 (.cout (\halfcarry[29] ), .sum (sum[30]), .cin (\halfcarry[28] )
    , .x (\halfsum[30] ), .y (\halfcout[29] ));
fullAdder__0_216 genblk2_28_f3 (.cout (\halfcarry[28] ), .sum (sum[29]), .cin (\halfcarry[27] )
    , .x (\halfsum[29] ), .y (\halfcout[28] ));
fullAdder__0_219 genblk2_27_f3 (.cout (\halfcarry[27] ), .sum (sum[28]), .cin (\halfcarry[26] )
    , .x (\halfsum[28] ), .y (\halfcout[27] ));
fullAdder__0_222 genblk2_26_f3 (.cout (\halfcarry[26] ), .sum (sum[27]), .cin (\halfcarry[25] )
    , .x (\halfsum[27] ), .y (\halfcout[26] ));
fullAdder__0_225 genblk2_25_f3 (.cout (\halfcarry[25] ), .sum (sum[26]), .cin (\halfcarry[24] )
    , .x (\halfsum[26] ), .y (\halfcout[25] ));
fullAdder__0_228 genblk2_24_f3 (.cout (\halfcarry[24] ), .sum (sum[25]), .cin (\halfcarry[23] )
    , .x (\halfsum[25] ), .y (\halfcout[24] ));
fullAdder__0_231 genblk2_23_f3 (.cout (\halfcarry[23] ), .sum (sum[24]), .cin (\halfcarry[22] )
    , .x (\halfsum[24] ), .y (\halfcout[23] ));
fullAdder__0_234 genblk2_22_f3 (.cout (\halfcarry[22] ), .sum (sum[23]), .cin (\halfcarry[21] )
    , .x (\halfsum[23] ), .y (\halfcout[22] ));
fullAdder__0_237 genblk2_21_f3 (.cout (\halfcarry[21] ), .sum (sum[22]), .cin (\halfcarry[20] )
    , .x (\halfsum[22] ), .y (\halfcout[21] ));
fullAdder__0_240 genblk2_20_f3 (.cout (\halfcarry[20] ), .sum (sum[21]), .cin (\halfcarry[19] )
    , .x (\halfsum[21] ), .y (\halfcout[20] ));
fullAdder__0_243 genblk2_19_f3 (.cout (\halfcarry[19] ), .sum (sum[20]), .cin (\halfcarry[18] )
    , .x (\halfsum[20] ), .y (\halfcout[19] ));
fullAdder__0_246 genblk2_18_f3 (.cout (\halfcarry[18] ), .sum (sum[19]), .cin (\halfcarry[17] )
    , .x (\halfsum[19] ), .y (\halfcout[18] ));
fullAdder__0_249 genblk2_17_f3 (.cout (\halfcarry[17] ), .sum (sum[18]), .cin (\halfcarry[16] )
    , .x (\halfsum[18] ), .y (\halfcout[17] ));
fullAdder__0_252 genblk2_16_f3 (.cout (\halfcarry[16] ), .sum (sum[17]), .cin (\halfcarry[15] )
    , .x (\halfsum[17] ), .y (\halfcout[16] ));
fullAdder__0_255 genblk2_15_f3 (.cout (\halfcarry[15] ), .sum (sum[16]), .cin (\halfcarry[14] )
    , .x (\halfsum[16] ), .y (\halfcout[15] ));
fullAdder__0_258 genblk2_14_f3 (.cout (\halfcarry[14] ), .sum (sum[15]), .cin (\halfcarry[13] )
    , .x (\halfsum[15] ), .y (\halfcout[14] ));
fullAdder__0_261 genblk2_13_f3 (.cout (\halfcarry[13] ), .sum (sum[14]), .cin (\halfcarry[12] )
    , .x (\halfsum[14] ), .y (\halfcout[13] ));
fullAdder__0_264 genblk2_12_f3 (.cout (\halfcarry[12] ), .sum (sum[13]), .cin (\halfcarry[11] )
    , .x (\halfsum[13] ), .y (\halfcout[12] ));
fullAdder__0_267 genblk2_11_f3 (.cout (\halfcarry[11] ), .sum (sum[12]), .cin (\halfcarry[10] )
    , .x (\halfsum[12] ), .y (\halfcout[11] ));
fullAdder__0_270 genblk2_10_f3 (.cout (\halfcarry[10] ), .sum (sum[11]), .cin (\halfcarry[9] )
    , .x (\halfsum[11] ), .y (\halfcout[10] ));
fullAdder__0_273 genblk2_9_f3 (.cout (\halfcarry[9] ), .sum (sum[10]), .cin (\halfcarry[8] )
    , .x (\halfsum[10] ), .y (\halfcout[9] ));
fullAdder__0_276 genblk2_8_f3 (.cout (\halfcarry[8] ), .sum (sum[9]), .cin (\halfcarry[7] )
    , .x (\halfsum[9] ), .y (\halfcout[8] ));
fullAdder__0_279 genblk2_7_f3 (.cout (\halfcarry[7] ), .sum (sum[8]), .cin (\halfcarry[6] )
    , .x (\halfsum[8] ), .y (\halfcout[7] ));
fullAdder__0_282 genblk2_6_f3 (.cout (\halfcarry[6] ), .sum (sum[7]), .cin (\halfcarry[5] )
    , .x (\halfsum[7] ), .y (\halfcout[6] ));
fullAdder__0_285 genblk2_5_f3 (.cout (\halfcarry[5] ), .sum (sum[6]), .cin (\halfcarry[4] )
    , .x (\halfsum[6] ), .y (\halfcout[5] ));
fullAdder__0_288 genblk2_4_f3 (.cout (\halfcarry[4] ), .sum (sum[5]), .cin (\halfcarry[3] )
    , .x (\halfsum[5] ), .y (\halfcout[4] ));
fullAdder__0_291 genblk2_3_f3 (.cout (\halfcarry[3] ), .sum (sum[4]), .cin (\halfcarry[2] )
    , .x (\halfsum[4] ), .y (\halfcout[3] ));
fullAdder__0_294 genblk2_2_f3 (.cout (\halfcarry[2] ), .sum (sum[3]), .cin (\halfcarry[1] )
    , .x (\halfsum[3] ), .y (\halfcout[2] ));
fullAdder__0_297 genblk2_1_f3 (.cout (\halfcarry[1] ), .sum (sum[2]), .cin (\halfcarry[0] )
    , .x (\halfsum[2] ), .y (\halfcout[1] ));
fullAdder__0_300 genblk1_31_fulladder_f1 (.sum (\halfsum[31] ), .x (a[31]), .y (b[31]));
fullAdder__0_303 genblk1_30_fulladder_f1 (.cout (\halfcout[30] ), .sum (\halfsum[30] )
    , .x (a[30]), .y (b[30]));
fullAdder__0_306 genblk1_29_fulladder_f1 (.cout (\halfcout[29] ), .sum (\halfsum[29] )
    , .x (a[29]), .y (b[29]));
fullAdder__0_309 genblk1_28_fulladder_f1 (.cout (\halfcout[28] ), .sum (\halfsum[28] )
    , .x (a[28]), .y (b[28]));
fullAdder__0_312 genblk1_27_fulladder_f1 (.cout (\halfcout[27] ), .sum (\halfsum[27] )
    , .x (a[27]), .y (b[27]));
fullAdder__0_315 genblk1_26_fulladder_f1 (.cout (\halfcout[26] ), .sum (\halfsum[26] )
    , .x (a[26]), .y (b[26]));
fullAdder__0_318 genblk1_25_fulladder_f1 (.cout (\halfcout[25] ), .sum (\halfsum[25] )
    , .x (a[25]), .y (b[25]));
fullAdder__0_321 genblk1_24_fulladder_f1 (.cout (\halfcout[24] ), .sum (\halfsum[24] )
    , .x (a[24]), .y (b[24]));
fullAdder__0_324 genblk1_23_fulladder_f1 (.cout (\halfcout[23] ), .sum (\halfsum[23] )
    , .x (a[23]), .y (b[23]));
fullAdder__0_327 genblk1_22_fulladder_f1 (.cout (\halfcout[22] ), .sum (\halfsum[22] )
    , .x (a[22]), .y (b[22]));
fullAdder__0_330 genblk1_21_fulladder_f1 (.cout (\halfcout[21] ), .sum (\halfsum[21] )
    , .x (a[21]), .y (b[21]));
fullAdder__0_333 genblk1_20_fulladder_f1 (.cout (\halfcout[20] ), .sum (\halfsum[20] )
    , .x (a[20]), .y (b[20]));
fullAdder__0_336 genblk1_19_fulladder_f1 (.cout (\halfcout[19] ), .sum (\halfsum[19] )
    , .x (a[19]), .y (b[19]));
fullAdder__0_339 genblk1_18_fulladder_f1 (.cout (\halfcout[18] ), .sum (\halfsum[18] )
    , .x (a[18]), .y (b[18]));
fullAdder__0_342 genblk1_17_fulladder_f1 (.cout (\halfcout[17] ), .sum (\halfsum[17] )
    , .x (a[17]), .y (b[17]));
fullAdder__0_345 genblk1_16_fulladder_f1 (.cout (\halfcout[16] ), .sum (\halfsum[16] )
    , .x (a[16]), .y (b[16]));
fullAdder__0_348 genblk1_15_fulladder_f1 (.cout (\halfcout[15] ), .sum (\halfsum[15] )
    , .x (a[15]), .y (b[15]));
fullAdder__0_351 genblk1_14_fulladder_f1 (.cout (\halfcout[14] ), .sum (\halfsum[14] )
    , .x (a[14]), .y (b[14]));
fullAdder__0_354 genblk1_13_fulladder_f1 (.cout (\halfcout[13] ), .sum (\halfsum[13] )
    , .x (a[13]), .y (b[13]));
fullAdder__0_357 genblk1_12_fulladder_f1 (.cout (\halfcout[12] ), .sum (\halfsum[12] )
    , .x (a[12]), .y (b[12]));
fullAdder__0_360 genblk1_11_fulladder_f1 (.cout (\halfcout[11] ), .sum (\halfsum[11] )
    , .x (a[11]), .y (b[11]));
fullAdder__0_363 genblk1_10_fulladder_f1 (.cout (\halfcout[10] ), .sum (\halfsum[10] )
    , .x (a[10]), .y (b[10]));
fullAdder__0_366 genblk1_9_fulladder_f1 (.cout (\halfcout[9] ), .sum (\halfsum[9] )
    , .x (a[9]), .y (b[9]));
fullAdder__0_369 genblk1_8_fulladder_f1 (.cout (\halfcout[8] ), .sum (\halfsum[8] )
    , .x (a[8]), .y (b[8]));
fullAdder__0_372 genblk1_7_fulladder_f1 (.cout (\halfcout[7] ), .sum (\halfsum[7] )
    , .x (a[7]), .y (b[7]));
fullAdder__0_375 genblk1_6_fulladder_f1 (.cout (\halfcout[6] ), .sum (\halfsum[6] )
    , .x (a[6]), .y (b[6]));
fullAdder__0_378 genblk1_5_fulladder_f1 (.cout (\halfcout[5] ), .sum (\halfsum[5] )
    , .x (a[5]), .y (b[5]));
fullAdder__0_381 genblk1_4_fulladder_f1 (.cout (\halfcout[4] ), .sum (\halfsum[4] )
    , .x (a[4]), .y (b[4]));
fullAdder__0_384 genblk1_3_fulladder_f1 (.cout (\halfcout[3] ), .sum (\halfsum[3] )
    , .x (a[3]), .y (b[3]));
fullAdder__0_387 genblk1_2_fulladder_f1 (.cout (\halfcout[2] ), .sum (\halfsum[2] )
    , .x (a[2]), .y (b[2]));
fullAdder__0_390 genblk1_1_fulladder_f1 (.cout (\halfcout[1] ), .sum (\halfsum[1] )
    , .x (a[1]), .y (b[1]));
fullAdder__0_393 genblk1_0_fulladder_f1 (.cout (\halfcout[0] ), .sum (sum[0]), .x (a[0]), .y (b[0]));
fullAdder__0_399 fulladder_f2 (.cout (\halfcarry[0] ), .sum (sum[1]), .x (\halfsum[1] ), .y (\halfcout[0] ));

endmodule //carrySaveAdder__0_400

module regFile__0_18 (clk_CTS_1_PP_0, clk_CTS_1_PP_1, read_data, read_data2, write_en, 
    write_data, write_data2, clk);

output [31:0] read_data2;
output [31:0] read_data;
output clk_CTS_1_PP_0;
input clk;
input [31:0] write_data2;
input [31:0] write_data;
input write_en;
input clk_CTS_1_PP_1;
wire CTS_n_tid0_2;
wire CTS_n_tid0_3;


CLKGATETST_X8 clk_gate_my_reg2_reg (.GCK (CTS_n_tid0_3), .CK (clk_CTS_1_PP_0), .E (write_en), .SE (1'b0 ));
DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid0_2), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid0_2), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid0_2), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid0_2), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid0_2), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid0_2), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid0_2), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid0_2), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid0_2), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid0_2), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid0_2), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid0_2), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid0_2), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid0_2), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid0_2), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid0_2), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid0_2), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid0_2), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid0_2), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid0_2), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid0_2), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid0_2), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid0_2), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid0_2), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid0_2), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid0_2), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid0_2), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid0_2), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid0_2), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid0_2), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid0_2), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid0_2), .D (write_data[31]));
DFF_X1 \my_reg2_reg[0]  (.Q (read_data2[0]), .CK (CTS_n_tid0_2), .D (write_data2[0]));
DFF_X1 \my_reg2_reg[1]  (.Q (read_data2[1]), .CK (CTS_n_tid0_2), .D (write_data2[1]));
DFF_X1 \my_reg2_reg[2]  (.Q (read_data2[2]), .CK (CTS_n_tid0_2), .D (write_data2[2]));
DFF_X1 \my_reg2_reg[3]  (.Q (read_data2[3]), .CK (CTS_n_tid0_2), .D (write_data2[3]));
DFF_X1 \my_reg2_reg[4]  (.Q (read_data2[4]), .CK (CTS_n_tid0_2), .D (write_data2[4]));
DFF_X1 \my_reg2_reg[5]  (.Q (read_data2[5]), .CK (CTS_n_tid0_2), .D (write_data2[5]));
DFF_X1 \my_reg2_reg[6]  (.Q (read_data2[6]), .CK (CTS_n_tid0_2), .D (write_data2[6]));
DFF_X1 \my_reg2_reg[7]  (.Q (read_data2[7]), .CK (CTS_n_tid0_2), .D (write_data2[7]));
DFF_X1 \my_reg2_reg[8]  (.Q (read_data2[8]), .CK (CTS_n_tid0_2), .D (write_data2[8]));
DFF_X1 \my_reg2_reg[9]  (.Q (read_data2[9]), .CK (CTS_n_tid0_2), .D (write_data2[9]));
DFF_X1 \my_reg2_reg[10]  (.Q (read_data2[10]), .CK (CTS_n_tid0_2), .D (write_data2[10]));
DFF_X1 \my_reg2_reg[11]  (.Q (read_data2[11]), .CK (CTS_n_tid0_2), .D (write_data2[11]));
DFF_X1 \my_reg2_reg[12]  (.Q (read_data2[12]), .CK (CTS_n_tid0_2), .D (write_data2[12]));
DFF_X1 \my_reg2_reg[13]  (.Q (read_data2[13]), .CK (CTS_n_tid0_2), .D (write_data2[13]));
DFF_X1 \my_reg2_reg[14]  (.Q (read_data2[14]), .CK (CTS_n_tid0_2), .D (write_data2[14]));
DFF_X1 \my_reg2_reg[15]  (.Q (read_data2[15]), .CK (CTS_n_tid0_2), .D (write_data2[15]));
DFF_X1 \my_reg2_reg[16]  (.Q (read_data2[16]), .CK (CTS_n_tid0_2), .D (write_data2[16]));
DFF_X1 \my_reg2_reg[17]  (.Q (read_data2[17]), .CK (CTS_n_tid0_2), .D (write_data2[17]));
DFF_X1 \my_reg2_reg[18]  (.Q (read_data2[18]), .CK (CTS_n_tid0_2), .D (write_data2[18]));
DFF_X1 \my_reg2_reg[19]  (.Q (read_data2[19]), .CK (CTS_n_tid0_2), .D (write_data2[19]));
DFF_X1 \my_reg2_reg[20]  (.Q (read_data2[20]), .CK (CTS_n_tid0_2), .D (write_data2[20]));
DFF_X1 \my_reg2_reg[21]  (.Q (read_data2[21]), .CK (CTS_n_tid0_2), .D (write_data2[21]));
DFF_X1 \my_reg2_reg[22]  (.Q (read_data2[22]), .CK (CTS_n_tid0_2), .D (write_data2[22]));
DFF_X1 \my_reg2_reg[23]  (.Q (read_data2[23]), .CK (CTS_n_tid0_2), .D (write_data2[23]));
DFF_X1 \my_reg2_reg[24]  (.Q (read_data2[24]), .CK (CTS_n_tid0_2), .D (write_data2[24]));
DFF_X1 \my_reg2_reg[25]  (.Q (read_data2[25]), .CK (CTS_n_tid0_2), .D (write_data2[25]));
DFF_X1 \my_reg2_reg[26]  (.Q (read_data2[26]), .CK (CTS_n_tid0_2), .D (write_data2[26]));
DFF_X1 \my_reg2_reg[27]  (.Q (read_data2[27]), .CK (CTS_n_tid0_2), .D (write_data2[27]));
DFF_X1 \my_reg2_reg[28]  (.Q (read_data2[28]), .CK (CTS_n_tid0_2), .D (write_data2[28]));
DFF_X1 \my_reg2_reg[29]  (.Q (read_data2[29]), .CK (CTS_n_tid0_2), .D (write_data2[29]));
DFF_X1 \my_reg2_reg[30]  (.Q (read_data2[30]), .CK (CTS_n_tid0_2), .D (write_data2[30]));
DFF_X1 \my_reg2_reg[31]  (.Q (read_data2[31]), .CK (CTS_n_tid0_2), .D (write_data2[31]));
CLKBUF_X3 CTS_L3_c_tid0_3 (.Z (CTS_n_tid0_2), .A (CTS_n_tid0_3));
CLKBUF_X2 CTS_L1_c_tid1_47 (.Z (clk_CTS_1_PP_0), .A (clk_CTS_1_PP_1));

endmodule //regFile__0_18

module BoothAlgo (M, Q, result, clk, start);

output [63:0] result;
input [31:0] M;
input [31:0] Q;
input clk;
input start;
wire CTS_n_tid1_147;
wire \read2[31] ;
wire \read2[30] ;
wire \read2[29] ;
wire \read2[28] ;
wire \read2[27] ;
wire \read2[26] ;
wire \read2[25] ;
wire \read2[24] ;
wire \read2[23] ;
wire \read2[22] ;
wire \read2[21] ;
wire \read2[20] ;
wire \read2[19] ;
wire \read2[18] ;
wire \read2[17] ;
wire \read2[16] ;
wire \read2[15] ;
wire \read2[14] ;
wire \read2[13] ;
wire \read2[12] ;
wire \read2[11] ;
wire \read2[10] ;
wire \read2[9] ;
wire \read2[8] ;
wire \read2[7] ;
wire \read2[6] ;
wire \read2[5] ;
wire \read2[4] ;
wire \read2[3] ;
wire \read2[2] ;
wire \read2[1] ;
wire \read2[0] ;
wire \read[31] ;
wire \read[30] ;
wire \read[29] ;
wire \read[28] ;
wire \read[27] ;
wire \read[26] ;
wire \read[25] ;
wire \read[24] ;
wire \read[23] ;
wire \read[22] ;
wire \read[21] ;
wire \read[20] ;
wire \read[19] ;
wire \read[18] ;
wire \read[17] ;
wire \read[16] ;
wire \read[15] ;
wire \read[14] ;
wire \read[13] ;
wire \read[12] ;
wire \read[11] ;
wire \read[10] ;
wire \read[9] ;
wire \read[8] ;
wire \read[7] ;
wire \read[6] ;
wire \read[5] ;
wire \read[4] ;
wire \read[3] ;
wire \read[2] ;
wire \read[1] ;
wire \read[0] ;
wire \SubM[31] ;
wire \SubM[30] ;
wire \SubM[29] ;
wire \SubM[28] ;
wire \SubM[27] ;
wire \SubM[26] ;
wire \SubM[25] ;
wire \SubM[24] ;
wire \SubM[23] ;
wire \SubM[22] ;
wire \SubM[21] ;
wire \SubM[20] ;
wire \SubM[19] ;
wire \SubM[18] ;
wire \SubM[17] ;
wire \SubM[16] ;
wire \SubM[15] ;
wire \SubM[14] ;
wire \SubM[13] ;
wire \SubM[12] ;
wire \SubM[11] ;
wire \SubM[10] ;
wire \SubM[9] ;
wire \SubM[8] ;
wire \SubM[7] ;
wire \SubM[6] ;
wire \SubM[5] ;
wire \SubM[4] ;
wire \SubM[3] ;
wire \SubM[2] ;
wire \SubM[1] ;
wire \SubM[0] ;
wire \AddM[31] ;
wire \AddM[30] ;
wire \AddM[29] ;
wire \AddM[28] ;
wire \AddM[27] ;
wire \AddM[26] ;
wire \AddM[25] ;
wire \AddM[24] ;
wire \AddM[23] ;
wire \AddM[22] ;
wire \AddM[21] ;
wire \AddM[20] ;
wire \AddM[19] ;
wire \AddM[18] ;
wire \AddM[17] ;
wire \AddM[16] ;
wire \AddM[15] ;
wire \AddM[14] ;
wire \AddM[13] ;
wire \AddM[12] ;
wire \AddM[11] ;
wire \AddM[10] ;
wire \AddM[9] ;
wire \AddM[8] ;
wire \AddM[7] ;
wire \AddM[6] ;
wire \AddM[5] ;
wire \AddM[4] ;
wire \AddM[3] ;
wire \AddM[2] ;
wire \AddM[1] ;
wire \AddM[0] ;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire \A[31] ;
wire \A[30] ;
wire \A[29] ;
wire \A[28] ;
wire \A[27] ;
wire \A[26] ;
wire \A[25] ;
wire \A[24] ;
wire \A[23] ;
wire \A[22] ;
wire \A[21] ;
wire \A[20] ;
wire \A[19] ;
wire \A[18] ;
wire \A[17] ;
wire \A[16] ;
wire \A[15] ;
wire \A[14] ;
wire \A[13] ;
wire \A[12] ;
wire \A[11] ;
wire \A[10] ;
wire \A[9] ;
wire \A[8] ;
wire \A[7] ;
wire \A[6] ;
wire \A[5] ;
wire \A[4] ;
wire \A[3] ;
wire \A[2] ;
wire \A[1] ;
wire \A[0] ;
wire n_0_102;
wire \l8[31] ;
wire \l8[30] ;
wire \l8[29] ;
wire \l8[28] ;
wire \l8[27] ;
wire \l8[26] ;
wire \l8[25] ;
wire \l8[24] ;
wire \l8[23] ;
wire \l8[22] ;
wire \l8[21] ;
wire \l8[20] ;
wire \l8[19] ;
wire \l8[18] ;
wire \l8[17] ;
wire \l8[16] ;
wire \l8[15] ;
wire \l8[14] ;
wire \l8[13] ;
wire \l8[12] ;
wire \l8[11] ;
wire \l8[10] ;
wire \l8[9] ;
wire \l8[8] ;
wire \l8[7] ;
wire \l8[6] ;
wire \l8[5] ;
wire \l8[4] ;
wire \l8[3] ;
wire \l8[2] ;
wire \l8[1] ;
wire \l8[0] ;
wire CTS_n_tid0_6;
wire \f8[31] ;
wire \f8[30] ;
wire \f8[29] ;
wire \f8[28] ;
wire \f8[27] ;
wire \f8[26] ;
wire \f8[25] ;
wire \f8[24] ;
wire \f8[23] ;
wire \f8[22] ;
wire \f8[21] ;
wire \f8[20] ;
wire \f8[19] ;
wire \f8[18] ;
wire \f8[17] ;
wire \f8[16] ;
wire \f8[15] ;
wire \f8[14] ;
wire \f8[13] ;
wire \f8[12] ;
wire \f8[11] ;
wire \f8[10] ;
wire \f8[9] ;
wire \f8[8] ;
wire \f8[7] ;
wire \f8[6] ;
wire \f8[5] ;
wire \f8[4] ;
wire \f8[3] ;
wire \f8[2] ;
wire \f8[1] ;
wire \f8[0] ;
wire write_en;
wire write_en2;
wire n_0_103;
wire \count[5] ;
wire \count[4] ;
wire \count[3] ;
wire \count[2] ;
wire \count[1] ;
wire \count[0] ;
wire q0;
wire CTS_n_tid1_7;
wire n_0_34;
wire n_0_35;
wire n_0_1_0;
wire n_0_36;
wire n_0_1_1;
wire n_0_37;
wire n_0_1_2;
wire n_0_38;
wire n_0_1_3;
wire n_0_39;
wire n_0_1_4;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_1_7;
wire n_0_40;
wire n_0_41;
wire n_0_1_8;
wire n_0_42;
wire n_0_1_9;
wire n_0_43;
wire n_0_1_10;
wire n_0_44;
wire n_0_1_11;
wire n_0_45;
wire n_0_1_12;
wire n_0_46;
wire n_0_1_13;
wire n_0_47;
wire n_0_1_14;
wire n_0_48;
wire n_0_1_15;
wire n_0_49;
wire n_0_1_16;
wire n_0_50;
wire n_0_1_17;
wire n_0_51;
wire n_0_1_18;
wire n_0_52;
wire n_0_1_19;
wire n_0_53;
wire n_0_1_20;
wire n_0_54;
wire n_0_1_21;
wire n_0_55;
wire n_0_1_22;
wire n_0_56;
wire n_0_1_23;
wire n_0_57;
wire n_0_1_24;
wire n_0_58;
wire n_0_1_25;
wire n_0_59;
wire n_0_1_26;
wire n_0_60;
wire n_0_1_27;
wire n_0_61;
wire n_0_1_28;
wire n_0_62;
wire n_0_1_29;
wire n_0_63;
wire n_0_1_30;
wire n_0_64;
wire n_0_1_31;
wire n_0_65;
wire n_0_1_32;
wire n_0_66;
wire n_0_1_33;
wire n_0_67;
wire n_0_1_34;
wire n_0_68;
wire n_0_1_35;
wire n_0_69;
wire n_0_1_36;
wire n_0_70;
wire n_0_1_37;
wire n_0_71;
wire n_0_1_38;
wire n_0_72;
wire n_0_1_39;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_1_40;
wire n_0_1_41;
wire n_0_1_42;
wire n_0_1_43;
wire n_0_101;
wire n_0_1_44;
wire n_0_1_45;
wire n_0_99;
wire n_0_100;
wire n_0_1_46;
wire n_0_1_47;
wire n_0_1_48;
wire n_0_33;
wire n_0_1_49;
wire uc_0;
wire drc_ipo_n3;
wire CTS_n_tid0_8;
wire CTS_n_tid1_9;
wire CTS_n_tid1_153;
wire CTS_n_tid1_154;
wire CTS_n_tid0_137;


INV_X1 i_0_1_124 (.ZN (n_0_1_49), .A (\l8[0] ));
INV_X1 i_0_1_123 (.ZN (n_0_33), .A (start));
NOR2_X1 i_0_1_122 (.ZN (n_0_1_48), .A1 (\count[1] ), .A2 (\count[0] ));
NAND2_X1 i_0_1_121 (.ZN (n_0_1_47), .A1 (\count[5] ), .A2 (n_0_1_48));
NOR4_X1 i_0_1_120 (.ZN (n_0_1_46), .A1 (n_0_1_47), .A2 (\count[2] ), .A3 (\count[3] ), .A4 (\count[4] ));
NAND2_X1 i_0_1_119 (.ZN (n_0_100), .A1 (n_0_1_46), .A2 (n_0_33));
NOR2_X1 i_0_1_118 (.ZN (n_0_99), .A1 (n_0_1_49), .A2 (start));
XNOR2_X1 i_0_1_117 (.ZN (n_0_1_45), .A (q0), .B (n_0_1_49));
NOR2_X4 i_0_1_116 (.ZN (n_0_1_44), .A1 (n_0_1_45), .A2 (start));
AOI21_X1 i_0_1_115 (.ZN (n_0_101), .A (n_0_1_44), .B1 (n_0_1_46), .B2 (n_0_33));
AND3_X2 i_0_1_114 (.ZN (n_0_1_43), .A1 (n_0_1_49), .A2 (n_0_33), .A3 (q0));
NOR3_X1 i_0_1_113 (.ZN (n_0_1_42), .A1 (n_0_1_49), .A2 (start), .A3 (q0));
AOI22_X1 i_0_1_112 (.ZN (n_0_1_41), .A1 (n_0_1_44), .A2 (\A[0] ), .B1 (start), .B2 (\read2[31] ));
AOI22_X1 i_0_1_111 (.ZN (n_0_1_40), .A1 (\AddM[0] ), .A2 (n_0_1_43), .B1 (drc_ipo_n3), .B2 (\SubM[0] ));
NAND2_X1 i_0_1_110 (.ZN (n_0_98), .A1 (n_0_1_41), .A2 (n_0_1_40));
MUX2_X1 i_0_1_109 (.Z (n_0_97), .A (\l8[31] ), .B (\read2[30] ), .S (start));
MUX2_X1 i_0_1_108 (.Z (n_0_96), .A (\l8[30] ), .B (\read2[29] ), .S (start));
MUX2_X1 i_0_1_107 (.Z (n_0_95), .A (\l8[29] ), .B (\read2[28] ), .S (start));
MUX2_X1 i_0_1_106 (.Z (n_0_94), .A (\l8[28] ), .B (\read2[27] ), .S (start));
MUX2_X1 i_0_1_105 (.Z (n_0_93), .A (\l8[27] ), .B (\read2[26] ), .S (start));
MUX2_X1 i_0_1_104 (.Z (n_0_92), .A (\l8[26] ), .B (\read2[25] ), .S (start));
MUX2_X1 i_0_1_103 (.Z (n_0_91), .A (\l8[25] ), .B (\read2[24] ), .S (start));
MUX2_X1 i_0_1_102 (.Z (n_0_90), .A (\l8[24] ), .B (\read2[23] ), .S (start));
MUX2_X1 i_0_1_101 (.Z (n_0_89), .A (\l8[23] ), .B (\read2[22] ), .S (start));
MUX2_X1 i_0_1_100 (.Z (n_0_88), .A (\l8[22] ), .B (\read2[21] ), .S (start));
MUX2_X1 i_0_1_99 (.Z (n_0_87), .A (\l8[21] ), .B (\read2[20] ), .S (start));
MUX2_X1 i_0_1_98 (.Z (n_0_86), .A (\l8[20] ), .B (\read2[19] ), .S (start));
MUX2_X1 i_0_1_97 (.Z (n_0_85), .A (\l8[19] ), .B (\read2[18] ), .S (start));
MUX2_X1 i_0_1_96 (.Z (n_0_84), .A (\l8[18] ), .B (\read2[17] ), .S (start));
MUX2_X1 i_0_1_95 (.Z (n_0_83), .A (\l8[17] ), .B (\read2[16] ), .S (start));
MUX2_X1 i_0_1_94 (.Z (n_0_82), .A (\l8[16] ), .B (\read2[15] ), .S (start));
MUX2_X1 i_0_1_93 (.Z (n_0_81), .A (\l8[15] ), .B (\read2[14] ), .S (start));
MUX2_X1 i_0_1_92 (.Z (n_0_80), .A (\l8[14] ), .B (\read2[13] ), .S (start));
MUX2_X1 i_0_1_91 (.Z (n_0_79), .A (\l8[13] ), .B (\read2[12] ), .S (start));
MUX2_X1 i_0_1_90 (.Z (n_0_78), .A (\l8[12] ), .B (\read2[11] ), .S (start));
MUX2_X1 i_0_1_89 (.Z (n_0_77), .A (\l8[11] ), .B (\read2[10] ), .S (start));
MUX2_X1 i_0_1_88 (.Z (n_0_76), .A (\l8[10] ), .B (\read2[9] ), .S (start));
MUX2_X1 i_0_1_87 (.Z (n_0_75), .A (\l8[9] ), .B (\read2[8] ), .S (start));
MUX2_X1 i_0_1_86 (.Z (n_0_74), .A (\l8[8] ), .B (\read2[7] ), .S (start));
MUX2_X1 i_0_1_85 (.Z (n_0_73), .A (\l8[7] ), .B (\read2[6] ), .S (start));
MUX2_X1 i_0_1_84 (.Z (n_0_109), .A (\l8[6] ), .B (\read2[5] ), .S (start));
MUX2_X1 i_0_1_83 (.Z (n_0_108), .A (\l8[5] ), .B (\read2[4] ), .S (start));
MUX2_X1 i_0_1_82 (.Z (n_0_107), .A (\l8[4] ), .B (\read2[3] ), .S (start));
MUX2_X1 i_0_1_81 (.Z (n_0_106), .A (\l8[3] ), .B (\read2[2] ), .S (start));
MUX2_X1 i_0_1_80 (.Z (n_0_105), .A (\l8[2] ), .B (\read2[1] ), .S (start));
MUX2_X1 i_0_1_79 (.Z (n_0_104), .A (\l8[1] ), .B (\read2[0] ), .S (start));
AOI22_X1 i_0_1_78 (.ZN (n_0_1_39), .A1 (\AddM[31] ), .A2 (n_0_1_43), .B1 (drc_ipo_n3), .B2 (\SubM[31] ));
INV_X1 i_0_1_77 (.ZN (n_0_72), .A (n_0_1_39));
NAND2_X1 i_0_1_76 (.ZN (n_0_1_38), .A1 (n_0_1_44), .A2 (\A[31] ));
NAND2_X1 i_0_1_75 (.ZN (n_0_71), .A1 (n_0_1_38), .A2 (n_0_1_39));
AOI222_X1 i_0_1_74 (.ZN (n_0_1_37), .A1 (n_0_1_44), .A2 (\A[30] ), .B1 (\SubM[30] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[30] ), .C2 (n_0_1_43));
INV_X1 i_0_1_73 (.ZN (n_0_70), .A (n_0_1_37));
AOI222_X1 i_0_1_72 (.ZN (n_0_1_36), .A1 (n_0_1_44), .A2 (\A[29] ), .B1 (\SubM[29] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[29] ), .C2 (n_0_1_43));
INV_X1 i_0_1_71 (.ZN (n_0_69), .A (n_0_1_36));
AOI222_X1 i_0_1_70 (.ZN (n_0_1_35), .A1 (n_0_1_44), .A2 (\A[28] ), .B1 (\SubM[28] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[28] ), .C2 (n_0_1_43));
INV_X1 i_0_1_69 (.ZN (n_0_68), .A (n_0_1_35));
AOI222_X1 i_0_1_68 (.ZN (n_0_1_34), .A1 (n_0_1_44), .A2 (\A[27] ), .B1 (\SubM[27] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[27] ), .C2 (n_0_1_43));
INV_X1 i_0_1_67 (.ZN (n_0_67), .A (n_0_1_34));
AOI222_X1 i_0_1_66 (.ZN (n_0_1_33), .A1 (n_0_1_44), .A2 (\A[26] ), .B1 (\SubM[26] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[26] ), .C2 (n_0_1_43));
INV_X1 i_0_1_65 (.ZN (n_0_66), .A (n_0_1_33));
AOI222_X1 i_0_1_64 (.ZN (n_0_1_32), .A1 (n_0_1_44), .A2 (\A[25] ), .B1 (\SubM[25] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[25] ), .C2 (n_0_1_43));
INV_X1 i_0_1_63 (.ZN (n_0_65), .A (n_0_1_32));
AOI222_X1 i_0_1_62 (.ZN (n_0_1_31), .A1 (n_0_1_44), .A2 (\A[24] ), .B1 (\SubM[24] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[24] ), .C2 (n_0_1_43));
INV_X1 i_0_1_61 (.ZN (n_0_64), .A (n_0_1_31));
AOI222_X1 i_0_1_60 (.ZN (n_0_1_30), .A1 (n_0_1_44), .A2 (\A[23] ), .B1 (\SubM[23] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[23] ), .C2 (n_0_1_43));
INV_X1 i_0_1_59 (.ZN (n_0_63), .A (n_0_1_30));
AOI222_X1 i_0_1_58 (.ZN (n_0_1_29), .A1 (n_0_1_44), .A2 (\A[22] ), .B1 (\SubM[22] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[22] ), .C2 (n_0_1_43));
INV_X1 i_0_1_57 (.ZN (n_0_62), .A (n_0_1_29));
AOI222_X1 i_0_1_56 (.ZN (n_0_1_28), .A1 (n_0_1_44), .A2 (\A[21] ), .B1 (\SubM[21] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[21] ), .C2 (n_0_1_43));
INV_X1 i_0_1_55 (.ZN (n_0_61), .A (n_0_1_28));
AOI222_X1 i_0_1_54 (.ZN (n_0_1_27), .A1 (n_0_1_44), .A2 (\A[20] ), .B1 (\SubM[20] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[20] ), .C2 (n_0_1_43));
INV_X1 i_0_1_53 (.ZN (n_0_60), .A (n_0_1_27));
AOI222_X1 i_0_1_52 (.ZN (n_0_1_26), .A1 (n_0_1_44), .A2 (\A[19] ), .B1 (\SubM[19] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[19] ), .C2 (n_0_1_43));
INV_X1 i_0_1_51 (.ZN (n_0_59), .A (n_0_1_26));
AOI222_X1 i_0_1_50 (.ZN (n_0_1_25), .A1 (n_0_1_44), .A2 (\A[18] ), .B1 (\SubM[18] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[18] ), .C2 (n_0_1_43));
INV_X1 i_0_1_49 (.ZN (n_0_58), .A (n_0_1_25));
AOI222_X1 i_0_1_48 (.ZN (n_0_1_24), .A1 (n_0_1_44), .A2 (\A[17] ), .B1 (\SubM[17] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[17] ), .C2 (n_0_1_43));
INV_X1 i_0_1_47 (.ZN (n_0_57), .A (n_0_1_24));
AOI222_X1 i_0_1_46 (.ZN (n_0_1_23), .A1 (n_0_1_44), .A2 (\A[16] ), .B1 (\SubM[16] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[16] ), .C2 (n_0_1_43));
INV_X1 i_0_1_45 (.ZN (n_0_56), .A (n_0_1_23));
AOI222_X1 i_0_1_44 (.ZN (n_0_1_22), .A1 (n_0_1_44), .A2 (\A[15] ), .B1 (\SubM[15] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[15] ), .C2 (n_0_1_43));
INV_X1 i_0_1_43 (.ZN (n_0_55), .A (n_0_1_22));
AOI222_X1 i_0_1_42 (.ZN (n_0_1_21), .A1 (n_0_1_44), .A2 (\A[14] ), .B1 (\SubM[14] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[14] ), .C2 (n_0_1_43));
INV_X1 i_0_1_41 (.ZN (n_0_54), .A (n_0_1_21));
AOI222_X1 i_0_1_40 (.ZN (n_0_1_20), .A1 (n_0_1_44), .A2 (\A[13] ), .B1 (\SubM[13] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[13] ), .C2 (n_0_1_43));
INV_X1 i_0_1_39 (.ZN (n_0_53), .A (n_0_1_20));
AOI222_X1 i_0_1_38 (.ZN (n_0_1_19), .A1 (n_0_1_44), .A2 (\A[12] ), .B1 (\SubM[12] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[12] ), .C2 (n_0_1_43));
INV_X1 i_0_1_37 (.ZN (n_0_52), .A (n_0_1_19));
AOI222_X1 i_0_1_36 (.ZN (n_0_1_18), .A1 (n_0_1_44), .A2 (\A[11] ), .B1 (\SubM[11] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[11] ), .C2 (n_0_1_43));
INV_X1 i_0_1_35 (.ZN (n_0_51), .A (n_0_1_18));
AOI222_X1 i_0_1_34 (.ZN (n_0_1_17), .A1 (n_0_1_44), .A2 (\A[10] ), .B1 (\SubM[10] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[10] ), .C2 (n_0_1_43));
INV_X1 i_0_1_33 (.ZN (n_0_50), .A (n_0_1_17));
AOI222_X1 i_0_1_32 (.ZN (n_0_1_16), .A1 (n_0_1_44), .A2 (\A[9] ), .B1 (\SubM[9] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[9] ), .C2 (n_0_1_43));
INV_X1 i_0_1_31 (.ZN (n_0_49), .A (n_0_1_16));
AOI222_X1 i_0_1_30 (.ZN (n_0_1_15), .A1 (n_0_1_44), .A2 (\A[8] ), .B1 (\SubM[8] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[8] ), .C2 (n_0_1_43));
INV_X1 i_0_1_29 (.ZN (n_0_48), .A (n_0_1_15));
AOI222_X1 i_0_1_28 (.ZN (n_0_1_14), .A1 (n_0_1_44), .A2 (\A[7] ), .B1 (\SubM[7] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[7] ), .C2 (n_0_1_43));
INV_X1 i_0_1_27 (.ZN (n_0_47), .A (n_0_1_14));
AOI222_X1 i_0_1_26 (.ZN (n_0_1_13), .A1 (n_0_1_44), .A2 (\A[6] ), .B1 (\SubM[6] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[6] ), .C2 (n_0_1_43));
INV_X1 i_0_1_25 (.ZN (n_0_46), .A (n_0_1_13));
AOI222_X1 i_0_1_24 (.ZN (n_0_1_12), .A1 (n_0_1_44), .A2 (\A[5] ), .B1 (\SubM[5] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[5] ), .C2 (n_0_1_43));
INV_X1 i_0_1_23 (.ZN (n_0_45), .A (n_0_1_12));
AOI222_X1 i_0_1_22 (.ZN (n_0_1_11), .A1 (n_0_1_44), .A2 (\A[4] ), .B1 (\SubM[4] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[4] ), .C2 (n_0_1_43));
INV_X1 i_0_1_21 (.ZN (n_0_44), .A (n_0_1_11));
AOI222_X1 i_0_1_20 (.ZN (n_0_1_10), .A1 (n_0_1_44), .A2 (\A[3] ), .B1 (\SubM[3] )
    , .B2 (drc_ipo_n3), .C1 (\AddM[3] ), .C2 (n_0_1_43));
INV_X1 i_0_1_19 (.ZN (n_0_43), .A (n_0_1_10));
AOI222_X1 i_0_1_18 (.ZN (n_0_1_9), .A1 (n_0_1_44), .A2 (\A[2] ), .B1 (\SubM[2] ), .B2 (drc_ipo_n3)
    , .C1 (\AddM[2] ), .C2 (n_0_1_43));
INV_X1 i_0_1_17 (.ZN (n_0_42), .A (n_0_1_9));
AOI222_X1 i_0_1_16 (.ZN (n_0_1_8), .A1 (n_0_1_44), .A2 (\A[1] ), .B1 (\SubM[1] ), .B2 (drc_ipo_n3)
    , .C1 (\AddM[1] ), .C2 (n_0_1_43));
INV_X1 i_0_1_15 (.ZN (n_0_41), .A (n_0_1_8));
OR2_X1 i_0_1_14 (.ZN (n_0_40), .A1 (start), .A2 (n_0_1_46));
AND3_X1 i_0_1_13 (.ZN (n_0_1_7), .A1 (\count[2] ), .A2 (\count[1] ), .A3 (\count[0] ));
AND2_X1 i_0_1_12 (.ZN (n_0_1_6), .A1 (\count[3] ), .A2 (n_0_1_7));
AND2_X1 i_0_1_11 (.ZN (n_0_1_5), .A1 (\count[4] ), .A2 (n_0_1_6));
XNOR2_X1 i_0_1_10 (.ZN (n_0_1_4), .A (\count[5] ), .B (n_0_1_5));
NOR2_X1 i_0_1_9 (.ZN (n_0_39), .A1 (start), .A2 (n_0_1_4));
OAI21_X1 i_0_1_8 (.ZN (n_0_1_3), .A (n_0_33), .B1 (\count[4] ), .B2 (n_0_1_6));
NOR2_X1 i_0_1_7 (.ZN (n_0_38), .A1 (n_0_1_5), .A2 (n_0_1_3));
OAI21_X1 i_0_1_6 (.ZN (n_0_1_2), .A (n_0_33), .B1 (\count[3] ), .B2 (n_0_1_7));
NOR2_X1 i_0_1_5 (.ZN (n_0_37), .A1 (n_0_1_6), .A2 (n_0_1_2));
AOI21_X1 i_0_1_4 (.ZN (n_0_1_1), .A (\count[2] ), .B1 (\count[1] ), .B2 (\count[0] ));
NOR3_X1 i_0_1_3 (.ZN (n_0_36), .A1 (start), .A2 (n_0_1_7), .A3 (n_0_1_1));
OAI21_X1 i_0_1_2 (.ZN (n_0_1_0), .A (n_0_33), .B1 (\count[1] ), .B2 (\count[0] ));
AOI21_X1 i_0_1_1 (.ZN (n_0_35), .A (n_0_1_0), .B1 (\count[0] ), .B2 (\count[1] ));
NOR2_X1 i_0_1_0 (.ZN (n_0_34), .A1 (start), .A2 (\count[0] ));
CLKGATETST_X8 clk_gate_A_reg__0 (.GCK (CTS_n_tid0_137), .CK (CTS_n_tid1_153), .E (n_0_100), .SE (1'b0 ));
DFF_X1 q0_reg (.Q (q0), .CK (CTS_n_tid0_6), .D (n_0_99));
DFF_X1 \count_reg[0]  (.Q (\count[0] ), .CK (CTS_n_tid0_6), .D (n_0_34));
DFF_X1 \count_reg[1]  (.Q (\count[1] ), .CK (CTS_n_tid0_8), .D (n_0_35));
DFF_X1 \count_reg[2]  (.Q (\count[2] ), .CK (CTS_n_tid0_8), .D (n_0_36));
DFF_X1 \count_reg[3]  (.Q (\count[3] ), .CK (CTS_n_tid0_6), .D (n_0_37));
DFF_X1 \count_reg[4]  (.Q (\count[4] ), .CK (CTS_n_tid0_8), .D (n_0_38));
DFF_X1 \count_reg[5]  (.Q (\count[5] ), .CK (CTS_n_tid0_8), .D (n_0_39));
MUX2_X1 write_en2_reg_enable_mux_0 (.Z (n_0_103), .A (write_en2), .B (n_0_33), .S (n_0_40));
DFF_X1 write_en2_reg (.Q (write_en2), .CK (CTS_n_tid1_147), .D (n_0_103));
DFF_X1 write_en_reg (.Q (write_en), .CK (CTS_n_tid1_147), .D (start));
DFF_X1 \f8_reg[0]  (.Q (\f8[0] ), .CK (CTS_n_tid1_7), .D (\read[0] ));
DFF_X1 \f8_reg[1]  (.Q (\f8[1] ), .CK (CTS_n_tid1_7), .D (\read[1] ));
DFF_X1 \f8_reg[2]  (.Q (\f8[2] ), .CK (CTS_n_tid1_7), .D (\read[2] ));
DFF_X1 \f8_reg[3]  (.Q (\f8[3] ), .CK (CTS_n_tid1_7), .D (\read[3] ));
DFF_X1 \f8_reg[4]  (.Q (\f8[4] ), .CK (CTS_n_tid1_7), .D (\read[4] ));
DFF_X1 \f8_reg[5]  (.Q (\f8[5] ), .CK (CTS_n_tid1_7), .D (\read[5] ));
DFF_X1 \f8_reg[6]  (.Q (\f8[6] ), .CK (CTS_n_tid1_7), .D (\read[6] ));
DFF_X1 \f8_reg[7]  (.Q (\f8[7] ), .CK (CTS_n_tid1_7), .D (\read[7] ));
DFF_X1 \f8_reg[8]  (.Q (\f8[8] ), .CK (CTS_n_tid1_7), .D (\read[8] ));
DFF_X1 \f8_reg[9]  (.Q (\f8[9] ), .CK (CTS_n_tid1_7), .D (\read[9] ));
DFF_X1 \f8_reg[10]  (.Q (\f8[10] ), .CK (CTS_n_tid1_7), .D (\read[10] ));
DFF_X1 \f8_reg[11]  (.Q (\f8[11] ), .CK (CTS_n_tid1_7), .D (\read[11] ));
DFF_X1 \f8_reg[12]  (.Q (\f8[12] ), .CK (CTS_n_tid1_7), .D (\read[12] ));
DFF_X1 \f8_reg[13]  (.Q (\f8[13] ), .CK (CTS_n_tid1_7), .D (\read[13] ));
DFF_X1 \f8_reg[14]  (.Q (\f8[14] ), .CK (CTS_n_tid1_7), .D (\read[14] ));
DFF_X1 \f8_reg[15]  (.Q (\f8[15] ), .CK (CTS_n_tid1_7), .D (\read[15] ));
DFF_X1 \f8_reg[16]  (.Q (\f8[16] ), .CK (CTS_n_tid1_7), .D (\read[16] ));
DFF_X1 \f8_reg[17]  (.Q (\f8[17] ), .CK (CTS_n_tid1_7), .D (\read[17] ));
DFF_X1 \f8_reg[18]  (.Q (\f8[18] ), .CK (CTS_n_tid1_7), .D (\read[18] ));
DFF_X1 \f8_reg[19]  (.Q (\f8[19] ), .CK (CTS_n_tid1_7), .D (\read[19] ));
DFF_X1 \f8_reg[20]  (.Q (\f8[20] ), .CK (CTS_n_tid1_7), .D (\read[20] ));
DFF_X1 \f8_reg[21]  (.Q (\f8[21] ), .CK (CTS_n_tid1_7), .D (\read[21] ));
DFF_X1 \f8_reg[22]  (.Q (\f8[22] ), .CK (CTS_n_tid1_7), .D (\read[22] ));
DFF_X1 \f8_reg[23]  (.Q (\f8[23] ), .CK (CTS_n_tid1_7), .D (\read[23] ));
DFF_X1 \f8_reg[24]  (.Q (\f8[24] ), .CK (CTS_n_tid1_7), .D (\read[24] ));
DFF_X1 \f8_reg[25]  (.Q (\f8[25] ), .CK (CTS_n_tid1_7), .D (\read[25] ));
DFF_X1 \f8_reg[26]  (.Q (\f8[26] ), .CK (CTS_n_tid1_7), .D (\read[26] ));
DFF_X1 \f8_reg[27]  (.Q (\f8[27] ), .CK (CTS_n_tid1_7), .D (\read[27] ));
DFF_X1 \f8_reg[28]  (.Q (\f8[28] ), .CK (CTS_n_tid1_7), .D (\read[28] ));
DFF_X1 \f8_reg[29]  (.Q (\f8[29] ), .CK (CTS_n_tid1_7), .D (\read[29] ));
DFF_X1 \f8_reg[30]  (.Q (\f8[30] ), .CK (CTS_n_tid1_7), .D (\read[30] ));
DFF_X1 \f8_reg[31]  (.Q (\f8[31] ), .CK (CTS_n_tid1_7), .D (\read[31] ));
CLKGATETST_X8 clk_gate_f8_reg (.GCK (CTS_n_tid1_9), .CK (CTS_n_tid1_153), .E (start), .SE (1'b0 ));
DFF_X1 \l8_reg[0]  (.Q (\l8[0] ), .CK (CTS_n_tid0_8), .D (n_0_104));
DFF_X1 \l8_reg[1]  (.Q (\l8[1] ), .CK (CTS_n_tid0_6), .D (n_0_105));
DFF_X1 \l8_reg[2]  (.Q (\l8[2] ), .CK (CTS_n_tid0_8), .D (n_0_106));
DFF_X1 \l8_reg[3]  (.Q (\l8[3] ), .CK (CTS_n_tid0_8), .D (n_0_107));
DFF_X1 \l8_reg[4]  (.Q (\l8[4] ), .CK (CTS_n_tid0_8), .D (n_0_108));
DFF_X1 \l8_reg[5]  (.Q (\l8[5] ), .CK (CTS_n_tid0_8), .D (n_0_109));
DFF_X1 \l8_reg[6]  (.Q (\l8[6] ), .CK (CTS_n_tid0_8), .D (n_0_73));
DFF_X1 \l8_reg[7]  (.Q (\l8[7] ), .CK (CTS_n_tid0_8), .D (n_0_74));
DFF_X1 \l8_reg[8]  (.Q (\l8[8] ), .CK (CTS_n_tid0_6), .D (n_0_75));
DFF_X1 \l8_reg[9]  (.Q (\l8[9] ), .CK (CTS_n_tid0_6), .D (n_0_76));
DFF_X1 \l8_reg[10]  (.Q (\l8[10] ), .CK (CTS_n_tid0_6), .D (n_0_77));
DFF_X1 \l8_reg[11]  (.Q (\l8[11] ), .CK (CTS_n_tid0_6), .D (n_0_78));
DFF_X1 \l8_reg[12]  (.Q (\l8[12] ), .CK (CTS_n_tid0_6), .D (n_0_79));
DFF_X1 \l8_reg[13]  (.Q (\l8[13] ), .CK (CTS_n_tid0_6), .D (n_0_80));
DFF_X1 \l8_reg[14]  (.Q (\l8[14] ), .CK (CTS_n_tid0_6), .D (n_0_81));
DFF_X1 \l8_reg[15]  (.Q (\l8[15] ), .CK (CTS_n_tid0_6), .D (n_0_82));
DFF_X1 \l8_reg[16]  (.Q (\l8[16] ), .CK (CTS_n_tid0_6), .D (n_0_83));
DFF_X1 \l8_reg[17]  (.Q (\l8[17] ), .CK (CTS_n_tid0_6), .D (n_0_84));
DFF_X1 \l8_reg[18]  (.Q (\l8[18] ), .CK (CTS_n_tid0_6), .D (n_0_85));
DFF_X1 \l8_reg[19]  (.Q (\l8[19] ), .CK (CTS_n_tid0_6), .D (n_0_86));
DFF_X1 \l8_reg[20]  (.Q (\l8[20] ), .CK (CTS_n_tid0_6), .D (n_0_87));
DFF_X1 \l8_reg[21]  (.Q (\l8[21] ), .CK (CTS_n_tid0_6), .D (n_0_88));
DFF_X1 \l8_reg[22]  (.Q (\l8[22] ), .CK (CTS_n_tid0_6), .D (n_0_89));
DFF_X1 \l8_reg[23]  (.Q (\l8[23] ), .CK (CTS_n_tid0_6), .D (n_0_90));
DFF_X1 \l8_reg[24]  (.Q (\l8[24] ), .CK (CTS_n_tid0_6), .D (n_0_91));
DFF_X1 \l8_reg[25]  (.Q (\l8[25] ), .CK (CTS_n_tid0_6), .D (n_0_92));
DFF_X1 \l8_reg[26]  (.Q (\l8[26] ), .CK (CTS_n_tid0_6), .D (n_0_93));
DFF_X1 \l8_reg[27]  (.Q (\l8[27] ), .CK (CTS_n_tid0_6), .D (n_0_94));
DFF_X1 \l8_reg[28]  (.Q (\l8[28] ), .CK (CTS_n_tid0_6), .D (n_0_95));
DFF_X1 \l8_reg[29]  (.Q (\l8[29] ), .CK (CTS_n_tid0_6), .D (n_0_96));
DFF_X1 \l8_reg[30]  (.Q (\l8[30] ), .CK (CTS_n_tid0_6), .D (n_0_97));
DFF_X1 \l8_reg[31]  (.Q (\l8[31] ), .CK (CTS_n_tid0_6), .D (n_0_98));
MUX2_X1 \A_reg[31]_enable_mux_0  (.Z (n_0_102), .A (\A[31] ), .B (n_0_72), .S (n_0_101));
DFF_X1 \A_reg[31]  (.Q (\A[31] ), .CK (CTS_n_tid1_147), .D (n_0_102));
DFF_X1 \A_reg[0]  (.Q (\A[0] ), .CK (CTS_n_tid0_6), .D (n_0_41));
DFF_X1 \A_reg[1]  (.Q (\A[1] ), .CK (CTS_n_tid0_6), .D (n_0_42));
DFF_X1 \A_reg[2]  (.Q (\A[2] ), .CK (CTS_n_tid0_6), .D (n_0_43));
DFF_X1 \A_reg[3]  (.Q (\A[3] ), .CK (CTS_n_tid0_6), .D (n_0_44));
DFF_X1 \A_reg[4]  (.Q (\A[4] ), .CK (CTS_n_tid0_6), .D (n_0_45));
DFF_X1 \A_reg[5]  (.Q (\A[5] ), .CK (CTS_n_tid0_6), .D (n_0_46));
DFF_X1 \A_reg[6]  (.Q (\A[6] ), .CK (CTS_n_tid0_6), .D (n_0_47));
DFF_X1 \A_reg[7]  (.Q (\A[7] ), .CK (CTS_n_tid0_6), .D (n_0_48));
DFF_X1 \A_reg[8]  (.Q (\A[8] ), .CK (CTS_n_tid0_6), .D (n_0_49));
DFF_X1 \A_reg[9]  (.Q (\A[9] ), .CK (CTS_n_tid0_8), .D (n_0_50));
DFF_X1 \A_reg[10]  (.Q (\A[10] ), .CK (CTS_n_tid0_6), .D (n_0_51));
DFF_X1 \A_reg[11]  (.Q (\A[11] ), .CK (CTS_n_tid0_8), .D (n_0_52));
DFF_X1 \A_reg[12]  (.Q (\A[12] ), .CK (CTS_n_tid0_8), .D (n_0_53));
DFF_X1 \A_reg[13]  (.Q (\A[13] ), .CK (CTS_n_tid0_8), .D (n_0_54));
DFF_X1 \A_reg[14]  (.Q (\A[14] ), .CK (CTS_n_tid0_8), .D (n_0_55));
DFF_X1 \A_reg[15]  (.Q (\A[15] ), .CK (CTS_n_tid0_8), .D (n_0_56));
DFF_X1 \A_reg[16]  (.Q (\A[16] ), .CK (CTS_n_tid0_8), .D (n_0_57));
DFF_X1 \A_reg[17]  (.Q (\A[17] ), .CK (CTS_n_tid0_8), .D (n_0_58));
DFF_X1 \A_reg[18]  (.Q (\A[18] ), .CK (CTS_n_tid0_8), .D (n_0_59));
DFF_X1 \A_reg[19]  (.Q (\A[19] ), .CK (CTS_n_tid0_8), .D (n_0_60));
DFF_X1 \A_reg[20]  (.Q (\A[20] ), .CK (CTS_n_tid0_8), .D (n_0_61));
DFF_X1 \A_reg[21]  (.Q (\A[21] ), .CK (CTS_n_tid0_8), .D (n_0_62));
DFF_X1 \A_reg[22]  (.Q (\A[22] ), .CK (CTS_n_tid0_8), .D (n_0_63));
DFF_X1 \A_reg[23]  (.Q (\A[23] ), .CK (CTS_n_tid0_8), .D (n_0_64));
DFF_X1 \A_reg[24]  (.Q (\A[24] ), .CK (CTS_n_tid0_8), .D (n_0_65));
DFF_X1 \A_reg[25]  (.Q (\A[25] ), .CK (CTS_n_tid0_8), .D (n_0_66));
DFF_X1 \A_reg[26]  (.Q (\A[26] ), .CK (CTS_n_tid0_8), .D (n_0_67));
DFF_X1 \A_reg[27]  (.Q (\A[27] ), .CK (CTS_n_tid0_8), .D (n_0_68));
DFF_X1 \A_reg[28]  (.Q (\A[28] ), .CK (CTS_n_tid0_8), .D (n_0_69));
DFF_X1 \A_reg[29]  (.Q (\A[29] ), .CK (CTS_n_tid0_8), .D (n_0_70));
DFF_X1 \A_reg[30]  (.Q (\A[30] ), .CK (CTS_n_tid0_8), .D (n_0_71));
datapath__0_17 i_0_0 (.p_0 ({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
    n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
    n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
    n_0_2, n_0_1, n_0_0, uc_0}), .f8 ({\f8[31] , \f8[30] , \f8[29] , \f8[28] , \f8[27] , 
    \f8[26] , \f8[25] , \f8[24] , \f8[23] , \f8[22] , \f8[21] , \f8[20] , \f8[19] , 
    \f8[18] , \f8[17] , \f8[16] , \f8[15] , \f8[14] , \f8[13] , \f8[12] , \f8[11] , 
    \f8[10] , \f8[9] , \f8[8] , \f8[7] , \f8[6] , \f8[5] , \f8[4] , \f8[3] , \f8[2] , 
    \f8[1] , \f8[0] }));
regFile inst2 (.read_data2 ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .read_data ({
    result[63], result[62], result[61], result[60], result[59], result[58], result[57], 
    result[56], result[55], result[54], result[53], result[52], result[51], result[50], 
    result[49], result[48], result[47], result[46], result[45], result[44], result[43], 
    result[42], result[41], result[40], result[39], result[38], result[37], result[36], 
    result[35], result[34], result[33], result[32]}), .write_data2 ({\l8[31] , \l8[30] , 
    \l8[29] , \l8[28] , \l8[27] , \l8[26] , \l8[25] , \l8[24] , \l8[23] , \l8[22] , 
    \l8[21] , \l8[20] , \l8[19] , \l8[18] , \l8[17] , \l8[16] , \l8[15] , \l8[14] , 
    \l8[13] , \l8[12] , \l8[11] , \l8[10] , \l8[9] , \l8[8] , \l8[7] , \l8[6] , \l8[5] , 
    \l8[4] , \l8[3] , \l8[2] , \l8[1] , \l8[0] }), .write_data ({\A[31] , \A[30] , 
    \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , 
    \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , 
    \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , 
    \A[1] , \A[0] }), .write_en (write_en2), .clk_CTS_1_PP_0 (CTS_n_tid1_154));
carrySaveAdder adder (.sum ({\AddM[31] , \AddM[30] , \AddM[29] , \AddM[28] , \AddM[27] , 
    \AddM[26] , \AddM[25] , \AddM[24] , \AddM[23] , \AddM[22] , \AddM[21] , \AddM[20] , 
    \AddM[19] , \AddM[18] , \AddM[17] , \AddM[16] , \AddM[15] , \AddM[14] , \AddM[13] , 
    \AddM[12] , \AddM[11] , \AddM[10] , \AddM[9] , \AddM[8] , \AddM[7] , \AddM[6] , 
    \AddM[5] , \AddM[4] , \AddM[3] , \AddM[2] , \AddM[1] , \AddM[0] }), .a ({\A[31] , 
    \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , 
    \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , 
    \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , 
    \A[2] , \A[1] , \A[0] }), .b ({\f8[31] , \f8[30] , \f8[29] , \f8[28] , \f8[27] , 
    \f8[26] , \f8[25] , \f8[24] , \f8[23] , \f8[22] , \f8[21] , \f8[20] , \f8[19] , 
    \f8[18] , \f8[17] , \f8[16] , \f8[15] , \f8[14] , \f8[13] , \f8[12] , \f8[11] , 
    \f8[10] , \f8[9] , \f8[8] , \f8[7] , \f8[6] , \f8[5] , \f8[4] , \f8[3] , \f8[2] , 
    \f8[1] , \f8[0] }));
carrySaveAdder__0_400 subtractor (.sum ({\SubM[31] , \SubM[30] , \SubM[29] , \SubM[28] , 
    \SubM[27] , \SubM[26] , \SubM[25] , \SubM[24] , \SubM[23] , \SubM[22] , \SubM[21] , 
    \SubM[20] , \SubM[19] , \SubM[18] , \SubM[17] , \SubM[16] , \SubM[15] , \SubM[14] , 
    \SubM[13] , \SubM[12] , \SubM[11] , \SubM[10] , \SubM[9] , \SubM[8] , \SubM[7] , 
    \SubM[6] , \SubM[5] , \SubM[4] , \SubM[3] , \SubM[2] , \SubM[1] , \SubM[0] })
    , .a ({\A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , 
    \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , 
    \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , 
    \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] }), .b ({n_0_30, n_0_29, n_0_28, 
    n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
    n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
    n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, \f8[0] }));
regFile__0_18 inst1 (.read_data2 ({\read2[31] , \read2[30] , \read2[29] , \read2[28] , 
    \read2[27] , \read2[26] , \read2[25] , \read2[24] , \read2[23] , \read2[22] , 
    \read2[21] , \read2[20] , \read2[19] , \read2[18] , \read2[17] , \read2[16] , 
    \read2[15] , \read2[14] , \read2[13] , \read2[12] , \read2[11] , \read2[10] , 
    \read2[9] , \read2[8] , \read2[7] , \read2[6] , \read2[5] , \read2[4] , \read2[3] , 
    \read2[2] , \read2[1] , \read2[0] }), .read_data ({\read[31] , \read[30] , \read[29] , 
    \read[28] , \read[27] , \read[26] , \read[25] , \read[24] , \read[23] , \read[22] , 
    \read[21] , \read[20] , \read[19] , \read[18] , \read[17] , \read[16] , \read[15] , 
    \read[14] , \read[13] , \read[12] , \read[11] , \read[10] , \read[9] , \read[8] , 
    \read[7] , \read[6] , \read[5] , \read[4] , \read[3] , \read[2] , \read[1] , 
    \read[0] }), .clk_CTS_1_PP_0 (CTS_n_tid1_154), .write_data2 ({Q[31], Q[30], Q[29], 
    Q[28], Q[27], Q[26], Q[25], Q[24], Q[23], Q[22], Q[21], Q[20], Q[19], Q[18], 
    Q[17], Q[16], Q[15], Q[14], Q[13], Q[12], Q[11], Q[10], Q[9], Q[8], Q[7], Q[6], 
    Q[5], Q[4], Q[3], Q[2], Q[1], Q[0]}), .write_data ({M[31], M[30], M[29], M[28], 
    M[27], M[26], M[25], M[24], M[23], M[22], M[21], M[20], M[19], M[18], M[17], 
    M[16], M[15], M[14], M[13], M[12], M[11], M[10], M[9], M[8], M[7], M[6], M[5], 
    M[4], M[3], M[2], M[1], M[0]}), .write_en (write_en), .clk_CTS_1_PP_1 (clk));
CLKBUF_X2 drc_ipo_c3 (.Z (drc_ipo_n3), .A (n_0_1_42));
CLKBUF_X3 CTS_L4_c_tid0_7 (.Z (CTS_n_tid0_6), .A (CTS_n_tid0_137));
CLKBUF_X3 CTS_L4_c_tid1_8 (.Z (CTS_n_tid1_7), .A (CTS_n_tid1_9));
CLKBUF_X3 CTS_L4_c_tid0_9 (.Z (CTS_n_tid0_8), .A (CTS_n_tid0_137));
CLKBUF_X1 CTS_L3_c_tid1_113 (.Z (CTS_n_tid1_147), .A (CTS_n_tid1_153));
CLKBUF_X2 CTS_L2_c_tid1_119 (.Z (CTS_n_tid1_153), .A (CTS_n_tid1_154));

endmodule //BoothAlgo


