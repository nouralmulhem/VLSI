/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 24 10:03:17 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 149233144 */

module regFile(read_data, read_data2, write_en, write_data, write_data2, clk);
   output [31:0]read_data;
   output [31:0]read_data2;
   input write_en;
   input [31:0]write_data;
   input [31:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[31]  (.D(write_data2[31]), .CK(n_0), .Q(read_data2[31]), 
      .QN());
   DFF_X1 \my_reg2_reg[30]  (.D(write_data2[30]), .CK(n_0), .Q(read_data2[30]), 
      .QN());
   DFF_X1 \my_reg2_reg[29]  (.D(write_data2[29]), .CK(n_0), .Q(read_data2[29]), 
      .QN());
   DFF_X1 \my_reg2_reg[28]  (.D(write_data2[28]), .CK(n_0), .Q(read_data2[28]), 
      .QN());
   DFF_X1 \my_reg2_reg[27]  (.D(write_data2[27]), .CK(n_0), .Q(read_data2[27]), 
      .QN());
   DFF_X1 \my_reg2_reg[26]  (.D(write_data2[26]), .CK(n_0), .Q(read_data2[26]), 
      .QN());
   DFF_X1 \my_reg2_reg[25]  (.D(write_data2[25]), .CK(n_0), .Q(read_data2[25]), 
      .QN());
   DFF_X1 \my_reg2_reg[24]  (.D(write_data2[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data2[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
   DFF_X1 \my_reg2_reg[22]  (.D(write_data2[22]), .CK(n_0), .Q(read_data2[22]), 
      .QN());
   DFF_X1 \my_reg2_reg[21]  (.D(write_data2[21]), .CK(n_0), .Q(read_data2[21]), 
      .QN());
   DFF_X1 \my_reg2_reg[20]  (.D(write_data2[20]), .CK(n_0), .Q(read_data2[20]), 
      .QN());
   DFF_X1 \my_reg2_reg[19]  (.D(write_data2[19]), .CK(n_0), .Q(read_data2[19]), 
      .QN());
   DFF_X1 \my_reg2_reg[18]  (.D(write_data2[18]), .CK(n_0), .Q(read_data2[18]), 
      .QN());
   DFF_X1 \my_reg2_reg[17]  (.D(write_data2[17]), .CK(n_0), .Q(read_data2[17]), 
      .QN());
   DFF_X1 \my_reg2_reg[16]  (.D(write_data2[16]), .CK(n_0), .Q(read_data2[16]), 
      .QN());
   DFF_X1 \my_reg2_reg[15]  (.D(write_data2[15]), .CK(n_0), .Q(read_data2[15]), 
      .QN());
   DFF_X1 \my_reg2_reg[14]  (.D(write_data2[14]), .CK(n_0), .Q(read_data2[14]), 
      .QN());
   DFF_X1 \my_reg2_reg[13]  (.D(write_data2[13]), .CK(n_0), .Q(read_data2[13]), 
      .QN());
   DFF_X1 \my_reg2_reg[12]  (.D(write_data2[12]), .CK(n_0), .Q(read_data2[12]), 
      .QN());
   DFF_X1 \my_reg2_reg[11]  (.D(write_data2[11]), .CK(n_0), .Q(read_data2[11]), 
      .QN());
   DFF_X1 \my_reg2_reg[10]  (.D(write_data2[10]), .CK(n_0), .Q(read_data2[10]), 
      .QN());
   DFF_X1 \my_reg2_reg[9]  (.D(write_data2[9]), .CK(n_0), .Q(read_data2[9]), 
      .QN());
   DFF_X1 \my_reg2_reg[8]  (.D(write_data2[8]), .CK(n_0), .Q(read_data2[8]), 
      .QN());
   DFF_X1 \my_reg2_reg[7]  (.D(write_data2[7]), .CK(n_0), .Q(read_data2[7]), 
      .QN());
   DFF_X1 \my_reg2_reg[6]  (.D(write_data2[6]), .CK(n_0), .Q(read_data2[6]), 
      .QN());
   DFF_X1 \my_reg2_reg[5]  (.D(write_data2[5]), .CK(n_0), .Q(read_data2[5]), 
      .QN());
   DFF_X1 \my_reg2_reg[4]  (.D(write_data2[4]), .CK(n_0), .Q(read_data2[4]), 
      .QN());
   DFF_X1 \my_reg2_reg[3]  (.D(write_data2[3]), .CK(n_0), .Q(read_data2[3]), 
      .QN());
   DFF_X1 \my_reg2_reg[2]  (.D(write_data2[2]), .CK(n_0), .Q(read_data2[2]), 
      .QN());
   DFF_X1 \my_reg2_reg[1]  (.D(write_data2[1]), .CK(n_0), .Q(read_data2[1]), 
      .QN());
   DFF_X1 \my_reg2_reg[0]  (.D(write_data2[0]), .CK(n_0), .Q(read_data2[0]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg2_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
endmodule

module full_adder__0_217(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
endmodule

module full_adder__0_221(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_225(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_229(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_233(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_237(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_241(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_245(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_249(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_253(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_257(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_261(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_265(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_269(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_273(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_277(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_281(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_285(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_289(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_293(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_297(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_301(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_305(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_309(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_313(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_317(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_321(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_325(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_329(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_333(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_337(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_341(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_345(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_349(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_353(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_357(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_361(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_365(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_369(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_373(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_377(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_381(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_385(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_389(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_393(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_397(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_401(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_405(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_409(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_413(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_417(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_421(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_425(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_429(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_433(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_437(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_441(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_445(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_449(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_453(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_457(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_461(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module full_adder__0_465(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_3), .ZN(o_sum));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_4), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(i_carry), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(i_carry), .A2(n_0_4), .ZN(n_0_3));
   XNOR2_X1 i_0_5 (.A(i_bit1), .B(i_bit2), .ZN(n_0_4));
endmodule

module full_adder(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_3), .ZN(o_sum));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_4), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(i_carry), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(i_carry), .A2(n_0_4), .ZN(n_0_3));
   XNOR2_X1 i_0_5 (.A(i_bit1), .B(i_bit2), .ZN(n_0_4));
endmodule

module carry_lookahead_adder(i_add1, i_add2, o_result, o_carry);
   input [63:0]i_add1;
   input [63:0]i_add2;
   output [63:0]o_result;
   output o_carry;

   wire n_0_38;
   wire n_0_21;
   wire n_0_27;
   wire n_0_39;
   wire n_0_40;
   wire n_0_35;
   wire n_0_41;
   wire n_0_42;
   wire w_G;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_155;
   wire n_0_157;
   wire n_0_47;
   wire n_0_167;
   wire n_0_168;
   wire n_0_48;
   wire n_0_201;
   wire n_0_202;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_237;
   wire n_0_49;
   wire n_0_259;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_50;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_51;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_181;
   wire n_0_389;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_171;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_146;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_111;
   wire n_0_19;
   wire n_0_101;
   wire n_0_20;
   wire n_0_22;
   wire n_0_96;
   wire n_0_23;
   wire n_0_223;
   wire n_0_219;
   wire n_0_216;
   wire n_0_235;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_209;
   wire n_0_213;
   wire n_0_238;
   wire n_0_191;
   wire n_0_186;
   wire n_0_28;
   wire n_0_29;
   wire n_0_176;
   wire n_0_30;
   wire n_0_166;
   wire n_0_161;
   wire n_0_151;
   wire n_0_31;
   wire n_0_32;
   wire n_0_141;
   wire n_0_131;
   wire n_0_126;
   wire n_0_33;
   wire n_0_121;
   wire n_0_34;
   wire n_0_116;
   wire n_0_36;
   wire n_0_37;
   wire n_0_106;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_156;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_169;
   wire n_0_170;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_214;
   wire n_0_215;
   wire n_0_217;
   wire n_0_218;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_234;
   wire n_0_236;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_260;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_296;
   wire n_0_297;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;

   full_adder__0_217 genblk1_0_full_adder_inst (.i_bit1(i_add1[0]), .i_bit2(
      i_add2[0]), .i_carry(), .o_sum(o_result[0]), .o_carry());
   full_adder__0_221 genblk1_1_full_adder_inst (.i_bit1(i_add1[1]), .i_bit2(
      i_add2[1]), .i_carry(w_G), .o_sum(o_result[1]), .o_carry());
   full_adder__0_225 genblk1_2_full_adder_inst (.i_bit1(i_add1[2]), .i_bit2(
      i_add2[2]), .i_carry(n_61), .o_sum(o_result[2]), .o_carry());
   full_adder__0_229 genblk1_3_full_adder_inst (.i_bit1(i_add1[3]), .i_bit2(
      i_add2[3]), .i_carry(n_23), .o_sum(o_result[3]), .o_carry());
   full_adder__0_233 genblk1_4_full_adder_inst (.i_bit1(i_add1[4]), .i_bit2(
      i_add2[4]), .i_carry(n_60), .o_sum(o_result[4]), .o_carry());
   full_adder__0_237 genblk1_5_full_adder_inst (.i_bit1(i_add1[5]), .i_bit2(
      i_add2[5]), .i_carry(n_22), .o_sum(o_result[5]), .o_carry());
   full_adder__0_241 genblk1_6_full_adder_inst (.i_bit1(i_add1[6]), .i_bit2(
      i_add2[6]), .i_carry(n_59), .o_sum(o_result[6]), .o_carry());
   full_adder__0_245 genblk1_7_full_adder_inst (.i_bit1(i_add1[7]), .i_bit2(
      i_add2[7]), .i_carry(n_21), .o_sum(o_result[7]), .o_carry());
   full_adder__0_249 genblk1_8_full_adder_inst (.i_bit1(i_add1[8]), .i_bit2(
      i_add2[8]), .i_carry(n_58), .o_sum(o_result[8]), .o_carry());
   full_adder__0_253 genblk1_9_full_adder_inst (.i_bit1(i_add1[9]), .i_bit2(
      i_add2[9]), .i_carry(n_57), .o_sum(o_result[9]), .o_carry());
   full_adder__0_257 genblk1_10_full_adder_inst (.i_bit1(i_add1[10]), .i_bit2(
      i_add2[10]), .i_carry(n_56), .o_sum(o_result[10]), .o_carry());
   full_adder__0_261 genblk1_11_full_adder_inst (.i_bit1(i_add1[11]), .i_bit2(
      i_add2[11]), .i_carry(n_20), .o_sum(o_result[11]), .o_carry());
   full_adder__0_265 genblk1_12_full_adder_inst (.i_bit1(i_add1[12]), .i_bit2(
      i_add2[12]), .i_carry(n_55), .o_sum(o_result[12]), .o_carry());
   full_adder__0_269 genblk1_13_full_adder_inst (.i_bit1(i_add1[13]), .i_bit2(
      i_add2[13]), .i_carry(n_19), .o_sum(o_result[13]), .o_carry());
   full_adder__0_273 genblk1_14_full_adder_inst (.i_bit1(i_add1[14]), .i_bit2(
      i_add2[14]), .i_carry(n_54), .o_sum(o_result[14]), .o_carry());
   full_adder__0_277 genblk1_15_full_adder_inst (.i_bit1(i_add1[15]), .i_bit2(
      i_add2[15]), .i_carry(n_18), .o_sum(o_result[15]), .o_carry());
   full_adder__0_281 genblk1_16_full_adder_inst (.i_bit1(i_add1[16]), .i_bit2(
      i_add2[16]), .i_carry(n_53), .o_sum(o_result[16]), .o_carry());
   full_adder__0_285 genblk1_17_full_adder_inst (.i_bit1(i_add1[17]), .i_bit2(
      i_add2[17]), .i_carry(n_52), .o_sum(o_result[17]), .o_carry());
   full_adder__0_289 genblk1_18_full_adder_inst (.i_bit1(i_add1[18]), .i_bit2(
      i_add2[18]), .i_carry(n_17), .o_sum(o_result[18]), .o_carry());
   full_adder__0_293 genblk1_19_full_adder_inst (.i_bit1(i_add1[19]), .i_bit2(
      i_add2[19]), .i_carry(n_24), .o_sum(o_result[19]), .o_carry());
   full_adder__0_297 genblk1_20_full_adder_inst (.i_bit1(i_add1[20]), .i_bit2(
      i_add2[20]), .i_carry(n_16), .o_sum(o_result[20]), .o_carry());
   full_adder__0_301 genblk1_21_full_adder_inst (.i_bit1(i_add1[21]), .i_bit2(
      i_add2[21]), .i_carry(n_25), .o_sum(o_result[21]), .o_carry());
   full_adder__0_305 genblk1_22_full_adder_inst (.i_bit1(i_add1[22]), .i_bit2(
      i_add2[22]), .i_carry(n_15), .o_sum(o_result[22]), .o_carry());
   full_adder__0_309 genblk1_23_full_adder_inst (.i_bit1(i_add1[23]), .i_bit2(
      i_add2[23]), .i_carry(n_26), .o_sum(o_result[23]), .o_carry());
   full_adder__0_313 genblk1_24_full_adder_inst (.i_bit1(i_add1[24]), .i_bit2(
      i_add2[24]), .i_carry(n_14), .o_sum(o_result[24]), .o_carry());
   full_adder__0_317 genblk1_25_full_adder_inst (.i_bit1(i_add1[25]), .i_bit2(
      i_add2[25]), .i_carry(n_27), .o_sum(o_result[25]), .o_carry());
   full_adder__0_321 genblk1_26_full_adder_inst (.i_bit1(i_add1[26]), .i_bit2(
      i_add2[26]), .i_carry(n_13), .o_sum(o_result[26]), .o_carry());
   full_adder__0_325 genblk1_27_full_adder_inst (.i_bit1(i_add1[27]), .i_bit2(
      i_add2[27]), .i_carry(n_28), .o_sum(o_result[27]), .o_carry());
   full_adder__0_329 genblk1_28_full_adder_inst (.i_bit1(i_add1[28]), .i_bit2(
      i_add2[28]), .i_carry(n_12), .o_sum(o_result[28]), .o_carry());
   full_adder__0_333 genblk1_29_full_adder_inst (.i_bit1(i_add1[29]), .i_bit2(
      i_add2[29]), .i_carry(n_29), .o_sum(o_result[29]), .o_carry());
   full_adder__0_337 genblk1_30_full_adder_inst (.i_bit1(i_add1[30]), .i_bit2(
      i_add2[30]), .i_carry(n_11), .o_sum(o_result[30]), .o_carry());
   full_adder__0_341 genblk1_31_full_adder_inst (.i_bit1(i_add1[31]), .i_bit2(
      i_add2[31]), .i_carry(n_30), .o_sum(o_result[31]), .o_carry());
   full_adder__0_345 genblk1_32_full_adder_inst (.i_bit1(i_add1[32]), .i_bit2(
      i_add2[32]), .i_carry(n_51), .o_sum(o_result[32]), .o_carry());
   full_adder__0_349 genblk1_33_full_adder_inst (.i_bit1(i_add1[33]), .i_bit2(
      i_add2[33]), .i_carry(n_31), .o_sum(o_result[33]), .o_carry());
   full_adder__0_353 genblk1_34_full_adder_inst (.i_bit1(i_add1[34]), .i_bit2(
      i_add2[34]), .i_carry(n_10), .o_sum(o_result[34]), .o_carry());
   full_adder__0_357 genblk1_35_full_adder_inst (.i_bit1(i_add1[35]), .i_bit2(
      i_add2[35]), .i_carry(n_32), .o_sum(o_result[35]), .o_carry());
   full_adder__0_361 genblk1_36_full_adder_inst (.i_bit1(i_add1[36]), .i_bit2(
      i_add2[36]), .i_carry(n_9), .o_sum(o_result[36]), .o_carry());
   full_adder__0_365 genblk1_37_full_adder_inst (.i_bit1(i_add1[37]), .i_bit2(
      i_add2[37]), .i_carry(n_33), .o_sum(o_result[37]), .o_carry());
   full_adder__0_369 genblk1_38_full_adder_inst (.i_bit1(i_add1[38]), .i_bit2(
      i_add2[38]), .i_carry(n_8), .o_sum(o_result[38]), .o_carry());
   full_adder__0_373 genblk1_39_full_adder_inst (.i_bit1(i_add1[39]), .i_bit2(
      i_add2[39]), .i_carry(n_34), .o_sum(o_result[39]), .o_carry());
   full_adder__0_377 genblk1_40_full_adder_inst (.i_bit1(i_add1[40]), .i_bit2(
      i_add2[40]), .i_carry(n_50), .o_sum(o_result[40]), .o_carry());
   full_adder__0_381 genblk1_41_full_adder_inst (.i_bit1(i_add1[41]), .i_bit2(
      i_add2[41]), .i_carry(n_35), .o_sum(o_result[41]), .o_carry());
   full_adder__0_385 genblk1_42_full_adder_inst (.i_bit1(i_add1[42]), .i_bit2(
      i_add2[42]), .i_carry(n_7), .o_sum(o_result[42]), .o_carry());
   full_adder__0_389 genblk1_43_full_adder_inst (.i_bit1(i_add1[43]), .i_bit2(
      i_add2[43]), .i_carry(n_36), .o_sum(o_result[43]), .o_carry());
   full_adder__0_393 genblk1_44_full_adder_inst (.i_bit1(i_add1[44]), .i_bit2(
      i_add2[44]), .i_carry(n_6), .o_sum(o_result[44]), .o_carry());
   full_adder__0_397 genblk1_45_full_adder_inst (.i_bit1(i_add1[45]), .i_bit2(
      i_add2[45]), .i_carry(n_37), .o_sum(o_result[45]), .o_carry());
   full_adder__0_401 genblk1_46_full_adder_inst (.i_bit1(i_add1[46]), .i_bit2(
      i_add2[46]), .i_carry(n_5), .o_sum(o_result[46]), .o_carry());
   full_adder__0_405 genblk1_47_full_adder_inst (.i_bit1(i_add1[47]), .i_bit2(
      i_add2[47]), .i_carry(n_38), .o_sum(o_result[47]), .o_carry());
   full_adder__0_409 genblk1_48_full_adder_inst (.i_bit1(i_add1[48]), .i_bit2(
      i_add2[48]), .i_carry(n_4), .o_sum(o_result[48]), .o_carry());
   full_adder__0_413 genblk1_49_full_adder_inst (.i_bit1(i_add1[49]), .i_bit2(
      i_add2[49]), .i_carry(n_39), .o_sum(o_result[49]), .o_carry());
   full_adder__0_417 genblk1_50_full_adder_inst (.i_bit1(i_add1[50]), .i_bit2(
      i_add2[50]), .i_carry(n_3), .o_sum(o_result[50]), .o_carry());
   full_adder__0_421 genblk1_51_full_adder_inst (.i_bit1(i_add1[51]), .i_bit2(
      i_add2[51]), .i_carry(n_40), .o_sum(o_result[51]), .o_carry());
   full_adder__0_425 genblk1_52_full_adder_inst (.i_bit1(i_add1[52]), .i_bit2(
      i_add2[52]), .i_carry(n_2), .o_sum(o_result[52]), .o_carry());
   full_adder__0_429 genblk1_53_full_adder_inst (.i_bit1(i_add1[53]), .i_bit2(
      i_add2[53]), .i_carry(n_41), .o_sum(o_result[53]), .o_carry());
   full_adder__0_433 genblk1_54_full_adder_inst (.i_bit1(i_add1[54]), .i_bit2(
      i_add2[54]), .i_carry(n_1), .o_sum(o_result[54]), .o_carry());
   full_adder__0_437 genblk1_55_full_adder_inst (.i_bit1(i_add1[55]), .i_bit2(
      i_add2[55]), .i_carry(n_44), .o_sum(o_result[55]), .o_carry());
   full_adder__0_441 genblk1_56_full_adder_inst (.i_bit1(i_add1[56]), .i_bit2(
      i_add2[56]), .i_carry(n_0), .o_sum(o_result[56]), .o_carry());
   full_adder__0_445 genblk1_57_full_adder_inst (.i_bit1(i_add1[57]), .i_bit2(
      i_add2[57]), .i_carry(n_42), .o_sum(o_result[57]), .o_carry());
   full_adder__0_449 genblk1_58_full_adder_inst (.i_bit1(i_add1[58]), .i_bit2(
      i_add2[58]), .i_carry(n_49), .o_sum(o_result[58]), .o_carry());
   full_adder__0_453 genblk1_59_full_adder_inst (.i_bit1(i_add1[59]), .i_bit2(
      i_add2[59]), .i_carry(n_45), .o_sum(o_result[59]), .o_carry());
   full_adder__0_457 genblk1_60_full_adder_inst (.i_bit1(i_add1[60]), .i_bit2(
      i_add2[60]), .i_carry(n_48), .o_sum(o_result[60]), .o_carry());
   full_adder__0_461 genblk1_61_full_adder_inst (.i_bit1(i_add1[61]), .i_bit2(
      i_add2[61]), .i_carry(n_43), .o_sum(o_result[61]), .o_carry());
   full_adder__0_465 genblk1_62_full_adder_inst (.i_bit1(i_add1[62]), .i_bit2(
      i_add2[62]), .i_carry(n_47), .o_sum(o_result[62]), .o_carry());
   full_adder genblk1_63_full_adder_inst (.i_bit1(i_add1[63]), .i_bit2(
      i_add2[63]), .i_carry(n_46), .o_sum(o_result[63]), .o_carry());
   INV_X1 i_0_0 (.A(n_0_96), .ZN(n_0));
   INV_X1 i_0_1 (.A(n_0_101), .ZN(n_1));
   INV_X1 i_0_2 (.A(n_0_106), .ZN(n_2));
   INV_X1 i_0_3 (.A(n_0_111), .ZN(n_3));
   INV_X1 i_0_4 (.A(n_0_116), .ZN(n_4));
   INV_X1 i_0_5 (.A(n_0_121), .ZN(n_5));
   OR2_X1 i_0_26 (.A1(i_add2[44]), .A2(i_add1[44]), .ZN(n_0_38));
   INV_X1 i_0_6 (.A(n_0_126), .ZN(n_6));
   INV_X1 i_0_7 (.A(n_0_131), .ZN(n_7));
   NAND2_X1 i_0_8 (.A1(i_add2[41]), .A2(i_add1[41]), .ZN(n_0_21));
   INV_X1 i_0_36 (.A(n_0_141), .ZN(n_8));
   INV_X1 i_0_9 (.A(n_0_146), .ZN(n_9));
   NAND2_X1 i_0_10 (.A1(i_add2[35]), .A2(i_add1[35]), .ZN(n_0_27));
   INV_X1 i_0_11 (.A(n_0_151), .ZN(n_10));
   OR2_X1 i_0_47 (.A1(i_add2[30]), .A2(i_add1[30]), .ZN(n_0_39));
   INV_X1 i_0_48 (.A(n_0_161), .ZN(n_11));
   NAND2_X1 i_0_49 (.A1(i_add2[29]), .A2(i_add1[29]), .ZN(n_0_40));
   INV_X1 i_0_12 (.A(n_0_166), .ZN(n_12));
   NAND2_X1 i_0_13 (.A1(i_add2[27]), .A2(i_add1[27]), .ZN(n_0_35));
   INV_X1 i_0_14 (.A(n_0_171), .ZN(n_13));
   INV_X1 i_0_15 (.A(n_0_176), .ZN(n_14));
   INV_X1 i_0_16 (.A(n_0_181), .ZN(n_15));
   NAND2_X1 i_0_17 (.A1(i_add2[21]), .A2(i_add1[21]), .ZN(n_0_41));
   INV_X1 i_0_18 (.A(n_0_186), .ZN(n_16));
   INV_X1 i_0_66 (.A(n_0_191), .ZN(n_17));
   NOR2_X1 i_0_71 (.A1(n_0_349), .A2(n_0_333), .ZN(n_18));
   NOR2_X1 i_0_74 (.A1(n_0_352), .A2(n_0_358), .ZN(n_19));
   NOR2_X1 i_0_77 (.A1(n_0_363), .A2(n_0_340), .ZN(n_20));
   NOR2_X1 i_0_19 (.A1(n_0_213), .A2(n_0_238), .ZN(n_21));
   NOR2_X1 i_0_89 (.A1(n_0_216), .A2(n_0_235), .ZN(n_22));
   OR2_X1 i_0_91 (.A1(i_add2[4]), .A2(i_add1[4]), .ZN(n_0_42));
   NOR2_X1 i_0_94 (.A1(n_0_223), .A2(n_0_219), .ZN(n_23));
   INV_X1 i_0_97 (.A(n_0_381), .ZN(w_G));
   BUF_X1 rt_shieldBuf__1 (.A(n_0_209), .Z(n_0_43));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(n_0_251), .Z(n_24));
   BUF_X1 rt_shieldBuf__1__1__1 (.A(n_0_28), .Z(n_25));
   BUF_X1 rt_shieldBuf__1__1__2 (.A(n_0_29), .Z(n_26));
   BUF_X1 rt_shieldBuf__1__1__3 (.A(n_0_30), .Z(n_27));
   BUF_X1 rt_shieldBuf__1__1__4 (.A(n_0_24), .Z(n_28));
   BUF_X1 rt_shieldBuf__1__1__5 (.A(n_0_233), .Z(n_29));
   BUF_X1 rt_shieldBuf__1__1__6 (.A(n_0_25), .Z(n_30));
   BUF_X1 rt_shieldBuf__1__1__7 (.A(n_0_261), .Z(n_31));
   BUF_X1 rt_shieldBuf__1__1__8 (.A(n_0_31), .Z(n_32));
   BUF_X1 rt_shieldBuf__1__1__9 (.A(n_0_32), .Z(n_33));
   BUF_X1 rt_shieldBuf__1__1__10 (.A(n_0_240), .Z(n_34));
   BUF_X1 rt_shieldBuf__1__1__11 (.A(n_0_26), .Z(n_35));
   BUF_X1 rt_shieldBuf__1__1__12 (.A(n_0_301), .Z(n_36));
   BUF_X1 rt_shieldBuf__1__1__13 (.A(n_0_33), .Z(n_37));
   BUF_X1 rt_shieldBuf__1__1__14 (.A(n_0_34), .Z(n_38));
   BUF_X1 rt_shieldBuf__1__1__15 (.A(n_0_36), .Z(n_39));
   BUF_X1 rt_shieldBuf__1__1__16 (.A(n_0_37), .Z(n_40));
   BUF_X1 rt_shieldBuf__1__1__17 (.A(n_0_52), .Z(n_41));
   INV_X1 i_0_159 (.A(n_0_369), .ZN(n_0_44));
   INV_X1 i_0_166 (.A(n_0_336), .ZN(n_0_45));
   INV_X1 i_0_176 (.A(n_0_178), .ZN(n_0_46));
   INV_X1 i_0_20 (.A(n_0_177), .ZN(n_0_155));
   OAI21_X1 i_0_21 (.A(n_0_255), .B1(n_0_256), .B2(n_0_155), .ZN(n_0_157));
   NAND2_X1 i_0_22 (.A1(n_0_157), .A2(n_0_175), .ZN(n_0_47));
   INV_X1 i_0_23 (.A(n_0_144), .ZN(n_0_167));
   NAND2_X1 i_0_24 (.A1(i_add1[20]), .A2(i_add2[20]), .ZN(n_0_168));
   OAI21_X1 i_0_188 (.A(n_0_41), .B1(n_0_167), .B2(n_0_168), .ZN(n_0_48));
   AND2_X1 i_0_25 (.A1(n_0_246), .A2(n_0_123), .ZN(n_0_201));
   INV_X1 i_0_27 (.A(n_0_122), .ZN(n_0_202));
   INV_X1 i_0_28 (.A(n_0_35), .ZN(n_0_230));
   OAI21_X1 i_0_29 (.A(n_0_119), .B1(n_0_201), .B2(n_0_230), .ZN(n_0_231));
   NAND2_X1 i_0_30 (.A1(i_add1[28]), .A2(i_add2[28]), .ZN(n_0_232));
   AOI21_X1 i_0_31 (.A(n_0_202), .B1(n_0_231), .B2(n_0_232), .ZN(n_0_233));
   OAI21_X1 i_0_32 (.A(n_0_232), .B1(n_0_35), .B2(n_0_120), .ZN(n_0_237));
   NAND2_X1 i_0_33 (.A1(n_0_237), .A2(n_0_122), .ZN(n_0_49));
   INV_X1 i_0_34 (.A(n_0_107), .ZN(n_0_259));
   AOI21_X1 i_0_35 (.A(n_0_259), .B1(n_0_326), .B2(n_0_156), .ZN(n_0_261));
   INV_X1 i_0_37 (.A(n_0_115), .ZN(n_0_262));
   NAND2_X1 i_0_38 (.A1(i_add1[34]), .A2(i_add2[34]), .ZN(n_0_263));
   OAI21_X1 i_0_39 (.A(n_0_27), .B1(n_0_262), .B2(n_0_263), .ZN(n_0_264));
   AOI22_X1 i_0_40 (.A1(n_0_264), .A2(n_0_113), .B1(i_add1[36]), .B2(i_add2[36]), 
      .ZN(n_0_50));
   AND3_X1 i_0_41 (.A1(n_0_124), .A2(n_0_84), .A3(n_0_99), .ZN(n_0_293));
   AND2_X1 i_0_42 (.A1(n_0_293), .A2(n_0_83), .ZN(n_0_294));
   INV_X1 i_0_43 (.A(n_0_82), .ZN(n_0_295));
   INV_X1 i_0_44 (.A(n_0_21), .ZN(n_0_298));
   OAI21_X1 i_0_45 (.A(n_0_80), .B1(n_0_294), .B2(n_0_298), .ZN(n_0_299));
   NAND2_X1 i_0_46 (.A1(i_add1[42]), .A2(i_add2[42]), .ZN(n_0_300));
   AOI21_X1 i_0_50 (.A(n_0_295), .B1(n_0_299), .B2(n_0_300), .ZN(n_0_301));
   OAI21_X1 i_0_51 (.A(n_0_300), .B1(n_0_21), .B2(n_0_81), .ZN(n_0_51));
   NOR3_X1 i_0_52 (.A1(n_0_195), .A2(n_0_184), .A3(n_0_174), .ZN(n_0_384));
   NOR2_X1 i_0_53 (.A1(n_0_384), .A2(n_0_147), .ZN(n_0_385));
   NAND2_X1 i_0_54 (.A1(n_0_385), .A2(n_0_143), .ZN(n_0_386));
   AOI21_X1 i_0_55 (.A(n_0_167), .B1(n_0_386), .B2(n_0_168), .ZN(n_0_387));
   INV_X1 i_0_56 (.A(n_0_41), .ZN(n_0_388));
   OAI21_X1 i_0_57 (.A(n_0_194), .B1(n_0_387), .B2(n_0_388), .ZN(n_0_181));
   NAND4_X1 i_0_58 (.A1(n_0_385), .A2(n_0_192), .A3(n_0_144), .A4(n_0_140), 
      .ZN(n_0_389));
   NAND2_X1 i_0_59 (.A1(n_0_389), .A2(n_0_189), .ZN(n_0_0));
   OAI22_X1 i_0_60 (.A1(n_0_0), .A2(n_0_183), .B1(i_add2[23]), .B2(i_add1[23]), 
      .ZN(n_0_1));
   INV_X1 i_0_61 (.A(n_0_138), .ZN(n_0_2));
   AOI21_X1 i_0_62 (.A(n_0_2), .B1(n_0_1), .B2(n_0_180), .ZN(n_0_3));
   INV_X1 i_0_63 (.A(n_0_139), .ZN(n_0_4));
   OAI21_X1 i_0_64 (.A(n_0_4), .B1(n_0_3), .B2(n_0_182), .ZN(n_0_171));
   NAND3_X1 i_0_65 (.A1(n_0_244), .A2(n_0_102), .A3(n_0_110), .ZN(n_0_5));
   AOI21_X1 i_0_67 (.A(n_0_262), .B1(n_0_5), .B2(n_0_263), .ZN(n_0_6));
   INV_X1 i_0_68 (.A(n_0_27), .ZN(n_0_7));
   OAI21_X1 i_0_69 (.A(n_0_113), .B1(n_0_6), .B2(n_0_7), .ZN(n_0_146));
   INV_X1 i_0_70 (.A(n_0_77), .ZN(n_0_8));
   AOI21_X1 i_0_72 (.A(n_0_66), .B1(n_0_293), .B2(n_0_8), .ZN(n_0_9));
   AOI21_X1 i_0_73 (.A(n_0_227), .B1(n_0_9), .B2(n_0_65), .ZN(n_0_10));
   INV_X1 i_0_75 (.A(n_0_97), .ZN(n_0_11));
   OAI21_X1 i_0_76 (.A(n_0_11), .B1(n_0_10), .B2(n_0_76), .ZN(n_0_12));
   INV_X1 i_0_78 (.A(n_0_98), .ZN(n_0_13));
   AOI21_X1 i_0_79 (.A(n_0_13), .B1(n_0_12), .B2(n_0_95), .ZN(n_0_14));
   INV_X1 i_0_80 (.A(n_0_94), .ZN(n_0_15));
   OAI21_X1 i_0_81 (.A(n_0_90), .B1(n_0_14), .B2(n_0_15), .ZN(n_0_16));
   AOI21_X1 i_0_82 (.A(n_0_93), .B1(n_0_16), .B2(n_0_63), .ZN(n_0_17));
   INV_X1 i_0_83 (.A(n_0_64), .ZN(n_0_18));
   OAI21_X1 i_0_84 (.A(n_0_91), .B1(n_0_17), .B2(n_0_18), .ZN(n_0_111));
   INV_X1 i_0_85 (.A(n_0_305), .ZN(n_0_19));
   OAI21_X1 i_0_86 (.A(n_0_286), .B1(n_0_52), .B2(n_0_19), .ZN(n_0_101));
   INV_X1 i_0_87 (.A(n_0_283), .ZN(n_0_20));
   AND3_X1 i_0_88 (.A1(n_0_297), .A2(n_0_292), .A3(n_0_20), .ZN(n_0_22));
   OAI21_X1 i_0_90 (.A(n_0_291), .B1(n_0_22), .B2(n_0_281), .ZN(n_0_96));
   NAND4_X1 i_0_92 (.A1(n_0_297), .A2(n_0_292), .A3(n_0_291), .A4(n_0_20), 
      .ZN(n_0_23));
   AOI21_X1 i_0_93 (.A(n_0_290), .B1(n_0_23), .B2(n_0_280), .ZN(n_42));
   BUF_X1 i_0_450 (.A(n_0_377), .Z(n_0_223));
   BUF_X1 i_0_451 (.A(n_0_376), .Z(n_0_219));
   BUF_X1 i_0_454 (.A(n_0_225), .Z(n_0_216));
   BUF_X1 i_0_455 (.A(n_0_234), .Z(n_0_235));
   BUF_X1 i_0_95 (.A(n_0_201), .Z(n_0_24));
   BUF_X1 i_0_96 (.A(n_0_328), .Z(n_0_25));
   BUF_X1 i_0_98 (.A(n_0_294), .Z(n_0_26));
   BUF_X1 i_0_464 (.A(n_0_319), .Z(n_43));
   BUF_X1 i_0_99 (.A(n_0_357), .Z(n_0_209));
   BUF_X1 i_0_100 (.A(n_0_367), .Z(n_0_213));
   BUF_X1 i_0_101 (.A(n_0_372), .Z(n_0_238));
   BUF_X1 i_0_472 (.A(n_0_252), .Z(n_0_191));
   BUF_X1 i_0_102 (.A(n_0_386), .Z(n_0_186));
   BUF_X1 i_0_103 (.A(n_0_387), .Z(n_0_28));
   BUF_X1 i_0_104 (.A(n_0_0), .Z(n_0_29));
   BUF_X1 i_0_105 (.A(n_0_1), .Z(n_0_176));
   BUF_X1 i_0_106 (.A(n_0_3), .Z(n_0_30));
   BUF_X1 i_0_107 (.A(n_0_231), .Z(n_0_166));
   BUF_X1 i_0_479 (.A(n_0_245), .Z(n_0_161));
   BUF_X1 i_0_108 (.A(n_0_5), .Z(n_0_151));
   BUF_X1 i_0_109 (.A(n_0_6), .Z(n_0_31));
   BUF_X1 i_0_482 (.A(n_0_242), .Z(n_0_32));
   BUF_X1 i_0_483 (.A(n_0_241), .Z(n_0_141));
   BUF_X1 i_0_110 (.A(n_0_299), .Z(n_0_131));
   BUF_X1 i_0_111 (.A(n_0_9), .Z(n_0_126));
   BUF_X1 i_0_112 (.A(n_0_10), .Z(n_0_33));
   BUF_X1 i_0_113 (.A(n_0_12), .Z(n_0_121));
   BUF_X1 i_0_114 (.A(n_0_14), .Z(n_0_34));
   BUF_X1 i_0_115 (.A(n_0_16), .Z(n_0_116));
   BUF_X1 i_0_116 (.A(n_0_17), .Z(n_0_36));
   BUF_X1 i_0_492 (.A(n_0_57), .Z(n_0_37));
   BUF_X1 i_0_117 (.A(n_0_54), .Z(n_0_106));
   BUF_X1 i_0_118 (.A(n_0_22), .Z(n_44));
   BUF_X1 i_0_496 (.A(n_0_323), .Z(n_45));
   AOI21_X1 i_0_119 (.A(n_0_226), .B1(n_0_54), .B2(n_0_53), .ZN(n_0_52));
   NAND2_X1 i_0_120 (.A1(i_add2[52]), .A2(i_add1[52]), .ZN(n_0_53));
   OAI22_X1 i_0_121 (.A1(i_add2[51]), .A2(i_add1[51]), .B1(n_0_57), .B2(n_0_55), 
      .ZN(n_0_54));
   INV_X1 i_0_122 (.A(n_0_56), .ZN(n_0_55));
   NAND2_X1 i_0_123 (.A1(i_add2[51]), .A2(i_add1[51]), .ZN(n_0_56));
   NAND2_X1 i_0_124 (.A1(n_0_68), .A2(n_0_59), .ZN(n_0_57));
   INV_X1 i_0_125 (.A(n_0_59), .ZN(n_0_58));
   AOI211_X1 i_0_126 (.A(n_0_61), .B(n_0_60), .C1(i_add2[50]), .C2(i_add1[50]), 
      .ZN(n_0_59));
   AOI211_X1 i_0_127 (.A(n_0_92), .B(n_0_72), .C1(n_0_64), .C2(n_0_63), .ZN(
      n_0_60));
   AOI21_X1 i_0_128 (.A(n_0_70), .B1(n_0_75), .B2(n_0_62), .ZN(n_0_61));
   AOI221_X1 i_0_129 (.A(n_0_66), .B1(i_add2[47]), .B2(i_add1[47]), .C1(
      i_add2[44]), .C2(i_add1[44]), .ZN(n_0_62));
   NAND2_X1 i_0_130 (.A1(i_add2[48]), .A2(i_add1[48]), .ZN(n_0_63));
   NAND2_X1 i_0_131 (.A1(i_add2[49]), .A2(i_add1[49]), .ZN(n_0_64));
   NAND2_X1 i_0_132 (.A1(i_add2[44]), .A2(i_add1[44]), .ZN(n_0_65));
   OAI22_X1 i_0_133 (.A1(n_0_239), .A2(n_0_236), .B1(n_0_79), .B2(n_0_67), 
      .ZN(n_0_66));
   NAND2_X1 i_0_134 (.A1(n_0_51), .A2(n_0_82), .ZN(n_0_67));
   NAND3_X1 i_0_135 (.A1(n_0_124), .A2(n_0_99), .A3(n_0_69), .ZN(n_0_68));
   NOR3_X1 i_0_136 (.A1(n_0_85), .A2(n_0_70), .A3(n_0_77), .ZN(n_0_69));
   NAND3_X1 i_0_137 (.A1(n_0_91), .A2(n_0_90), .A3(n_0_71), .ZN(n_0_70));
   AOI211_X1 i_0_138 (.A(n_0_93), .B(n_0_72), .C1(n_0_94), .C2(n_0_73), .ZN(
      n_0_71));
   NOR2_X1 i_0_139 (.A1(i_add2[50]), .A2(i_add1[50]), .ZN(n_0_72));
   NAND2_X1 i_0_140 (.A1(n_0_98), .A2(n_0_74), .ZN(n_0_73));
   OAI21_X1 i_0_141 (.A(n_0_75), .B1(n_0_227), .B2(n_0_97), .ZN(n_0_74));
   AOI21_X1 i_0_142 (.A(n_0_76), .B1(i_add2[46]), .B2(i_add1[46]), .ZN(n_0_75));
   AND2_X1 i_0_143 (.A1(i_add2[45]), .A2(i_add1[45]), .ZN(n_0_76));
   NAND4_X1 i_0_144 (.A1(n_0_83), .A2(n_0_82), .A3(n_0_80), .A4(n_0_78), 
      .ZN(n_0_77));
   INV_X1 i_0_145 (.A(n_0_79), .ZN(n_0_78));
   NOR2_X1 i_0_146 (.A1(i_add2[43]), .A2(i_add1[43]), .ZN(n_0_79));
   INV_X1 i_0_147 (.A(n_0_81), .ZN(n_0_80));
   NOR2_X1 i_0_148 (.A1(i_add2[41]), .A2(i_add1[41]), .ZN(n_0_81));
   OR2_X1 i_0_149 (.A1(i_add2[42]), .A2(i_add1[42]), .ZN(n_0_82));
   OR2_X1 i_0_150 (.A1(i_add2[40]), .A2(i_add1[40]), .ZN(n_0_83));
   INV_X1 i_0_151 (.A(n_0_85), .ZN(n_0_84));
   AOI21_X1 i_0_152 (.A(n_0_86), .B1(i_add2[40]), .B2(i_add1[40]), .ZN(n_0_85));
   AOI21_X1 i_0_153 (.A(n_0_88), .B1(n_0_128), .B2(n_0_87), .ZN(n_0_86));
   OAI21_X1 i_0_154 (.A(n_0_89), .B1(i_add2[37]), .B2(i_add1[37]), .ZN(n_0_87));
   NOR2_X1 i_0_155 (.A1(i_add2[39]), .A2(i_add1[39]), .ZN(n_0_88));
   OR2_X1 i_0_156 (.A1(i_add2[38]), .A2(i_add1[38]), .ZN(n_0_89));
   OR2_X1 i_0_157 (.A1(i_add2[47]), .A2(i_add1[47]), .ZN(n_0_90));
   INV_X1 i_0_158 (.A(n_0_92), .ZN(n_0_91));
   NOR2_X1 i_0_160 (.A1(i_add2[49]), .A2(i_add1[49]), .ZN(n_0_92));
   NOR2_X1 i_0_161 (.A1(i_add2[48]), .A2(i_add1[48]), .ZN(n_0_93));
   NAND2_X1 i_0_162 (.A1(i_add2[47]), .A2(i_add1[47]), .ZN(n_0_94));
   NAND2_X1 i_0_163 (.A1(i_add2[46]), .A2(i_add1[46]), .ZN(n_0_95));
   NOR2_X1 i_0_164 (.A1(i_add2[45]), .A2(i_add1[45]), .ZN(n_0_97));
   OR2_X1 i_0_165 (.A1(i_add2[46]), .A2(i_add1[46]), .ZN(n_0_98));
   NAND2_X1 i_0_167 (.A1(n_0_125), .A2(n_0_100), .ZN(n_0_99));
   OAI211_X1 i_0_168 (.A(n_0_108), .B(n_0_102), .C1(n_0_130), .C2(n_0_117), 
      .ZN(n_0_100));
   NAND2_X1 i_0_169 (.A1(n_0_153), .A2(n_0_103), .ZN(n_0_102));
   NAND2_X1 i_0_170 (.A1(n_0_107), .A2(n_0_104), .ZN(n_0_103));
   OAI21_X1 i_0_171 (.A(n_0_154), .B1(n_0_228), .B2(n_0_105), .ZN(n_0_104));
   NOR2_X1 i_0_172 (.A1(i_add2[31]), .A2(i_add1[31]), .ZN(n_0_105));
   OR2_X1 i_0_173 (.A1(i_add2[32]), .A2(i_add1[32]), .ZN(n_0_107));
   NOR3_X1 i_0_174 (.A1(n_0_114), .A2(n_0_109), .A3(n_0_112), .ZN(n_0_108));
   OAI21_X1 i_0_175 (.A(n_0_115), .B1(i_add2[36]), .B2(i_add1[36]), .ZN(n_0_109));
   INV_X1 i_0_177 (.A(n_0_112), .ZN(n_0_110));
   NOR2_X1 i_0_178 (.A1(i_add2[33]), .A2(i_add1[33]), .ZN(n_0_112));
   INV_X1 i_0_179 (.A(n_0_114), .ZN(n_0_113));
   NOR2_X1 i_0_180 (.A1(i_add2[35]), .A2(i_add1[35]), .ZN(n_0_114));
   OR2_X1 i_0_181 (.A1(i_add2[34]), .A2(i_add1[34]), .ZN(n_0_115));
   INV_X1 i_0_182 (.A(n_0_118), .ZN(n_0_117));
   NAND4_X1 i_0_183 (.A1(n_0_123), .A2(n_0_122), .A3(n_0_119), .A4(n_0_162), 
      .ZN(n_0_118));
   INV_X1 i_0_184 (.A(n_0_120), .ZN(n_0_119));
   NOR2_X1 i_0_185 (.A1(i_add2[27]), .A2(i_add1[27]), .ZN(n_0_120));
   OR2_X1 i_0_186 (.A1(i_add2[28]), .A2(i_add1[28]), .ZN(n_0_122));
   OR2_X1 i_0_187 (.A1(i_add2[26]), .A2(i_add1[26]), .ZN(n_0_123));
   OAI211_X1 i_0_189 (.A(n_0_132), .B(n_0_125), .C1(n_0_134), .C2(n_0_133), 
      .ZN(n_0_124));
   AND4_X1 i_0_190 (.A1(n_0_149), .A2(n_0_127), .A3(n_0_164), .A4(n_0_128), 
      .ZN(n_0_125));
   NAND2_X1 i_0_191 (.A1(i_add2[40]), .A2(i_add1[40]), .ZN(n_0_127));
   AOI21_X1 i_0_192 (.A(n_0_129), .B1(i_add2[38]), .B2(i_add1[38]), .ZN(n_0_128));
   AND2_X1 i_0_193 (.A1(i_add2[39]), .A2(i_add1[39]), .ZN(n_0_129));
   INV_X1 i_0_194 (.A(n_0_132), .ZN(n_0_130));
   NOR2_X1 i_0_195 (.A1(n_0_160), .A2(n_0_152), .ZN(n_0_132));
   NOR2_X1 i_0_196 (.A1(n_0_195), .A2(n_0_165), .ZN(n_0_133));
   OAI22_X1 i_0_197 (.A1(n_0_169), .A2(n_0_137), .B1(n_0_173), .B2(n_0_135), 
      .ZN(n_0_134));
   AOI21_X1 i_0_198 (.A(n_0_139), .B1(n_0_170), .B2(n_0_136), .ZN(n_0_135));
   OAI21_X1 i_0_199 (.A(n_0_138), .B1(i_add2[23]), .B2(i_add1[23]), .ZN(n_0_136));
   NOR4_X1 i_0_200 (.A1(n_0_147), .A2(n_0_145), .A3(n_0_142), .A4(n_0_193), 
      .ZN(n_0_137));
   OR2_X1 i_0_201 (.A1(i_add2[24]), .A2(i_add1[24]), .ZN(n_0_138));
   NOR2_X1 i_0_202 (.A1(i_add2[25]), .A2(i_add1[25]), .ZN(n_0_139));
   INV_X1 i_0_203 (.A(n_0_142), .ZN(n_0_140));
   NAND2_X1 i_0_204 (.A1(n_0_194), .A2(n_0_143), .ZN(n_0_142));
   OR2_X1 i_0_205 (.A1(i_add2[19]), .A2(i_add1[19]), .ZN(n_0_143));
   INV_X1 i_0_206 (.A(n_0_145), .ZN(n_0_144));
   NOR2_X1 i_0_207 (.A1(i_add2[20]), .A2(i_add1[20]), .ZN(n_0_145));
   AOI21_X1 i_0_208 (.A(n_0_46), .B1(n_0_47), .B2(n_0_258), .ZN(n_0_147));
   NAND2_X1 i_0_209 (.A1(i_add2[38]), .A2(i_add1[38]), .ZN(n_0_148));
   NAND2_X1 i_0_210 (.A1(i_add2[37]), .A2(i_add1[37]), .ZN(n_0_149));
   INV_X1 i_0_211 (.A(n_0_152), .ZN(n_0_150));
   NAND3_X1 i_0_212 (.A1(n_0_158), .A2(n_0_153), .A3(n_0_154), .ZN(n_0_152));
   NAND2_X1 i_0_213 (.A1(i_add2[33]), .A2(i_add1[33]), .ZN(n_0_153));
   AND2_X1 i_0_214 (.A1(n_0_159), .A2(n_0_156), .ZN(n_0_154));
   NAND2_X1 i_0_215 (.A1(i_add2[32]), .A2(i_add1[32]), .ZN(n_0_156));
   NAND2_X1 i_0_216 (.A1(i_add2[30]), .A2(i_add1[30]), .ZN(n_0_158));
   NAND2_X1 i_0_217 (.A1(i_add2[31]), .A2(i_add1[31]), .ZN(n_0_159));
   AOI21_X1 i_0_218 (.A(n_0_163), .B1(n_0_49), .B2(n_0_40), .ZN(n_0_160));
   INV_X1 i_0_219 (.A(n_0_163), .ZN(n_0_162));
   NOR2_X1 i_0_220 (.A1(i_add2[29]), .A2(i_add1[29]), .ZN(n_0_163));
   OAI21_X1 i_0_221 (.A(n_0_229), .B1(i_add2[36]), .B2(i_add1[36]), .ZN(n_0_164));
   OR3_X1 i_0_222 (.A1(n_0_184), .A2(n_0_174), .A3(n_0_169), .ZN(n_0_165));
   NAND3_X1 i_0_223 (.A1(n_0_172), .A2(n_0_170), .A3(n_0_189), .ZN(n_0_169));
   AOI21_X1 i_0_224 (.A(n_0_182), .B1(i_add2[24]), .B2(i_add1[24]), .ZN(n_0_170));
   NOR2_X1 i_0_225 (.A1(n_0_183), .A2(n_0_173), .ZN(n_0_172));
   AND2_X1 i_0_226 (.A1(i_add2[26]), .A2(i_add1[26]), .ZN(n_0_173));
   NAND4_X1 i_0_227 (.A1(n_0_179), .A2(n_0_178), .A3(n_0_177), .A4(n_0_175), 
      .ZN(n_0_174));
   NAND2_X1 i_0_228 (.A1(i_add2[18]), .A2(i_add1[18]), .ZN(n_0_175));
   NAND2_X1 i_0_229 (.A1(i_add2[17]), .A2(i_add1[17]), .ZN(n_0_177));
   NAND2_X1 i_0_230 (.A1(i_add2[19]), .A2(i_add1[19]), .ZN(n_0_178));
   NAND2_X1 i_0_231 (.A1(i_add2[16]), .A2(i_add1[16]), .ZN(n_0_179));
   NAND2_X1 i_0_232 (.A1(i_add2[24]), .A2(i_add1[24]), .ZN(n_0_180));
   AND2_X1 i_0_233 (.A1(i_add2[25]), .A2(i_add1[25]), .ZN(n_0_182));
   AND2_X1 i_0_234 (.A1(i_add2[23]), .A2(i_add1[23]), .ZN(n_0_183));
   OAI21_X1 i_0_235 (.A(n_0_187), .B1(n_0_188), .B2(n_0_185), .ZN(n_0_184));
   OAI21_X1 i_0_236 (.A(n_0_332), .B1(n_0_344), .B2(n_0_45), .ZN(n_0_185));
   NAND2_X1 i_0_237 (.A1(i_add2[15]), .A2(i_add1[15]), .ZN(n_0_187));
   NOR2_X1 i_0_238 (.A1(i_add2[15]), .A2(i_add1[15]), .ZN(n_0_188));
   AOI22_X1 i_0_239 (.A1(i_add2[22]), .A2(i_add1[22]), .B1(n_0_192), .B2(n_0_190), 
      .ZN(n_0_189));
   AND2_X1 i_0_240 (.A1(n_0_48), .A2(n_0_194), .ZN(n_0_190));
   INV_X1 i_0_241 (.A(n_0_193), .ZN(n_0_192));
   NOR2_X1 i_0_242 (.A1(i_add2[22]), .A2(i_add1[22]), .ZN(n_0_193));
   OR2_X1 i_0_243 (.A1(i_add2[21]), .A2(i_add1[21]), .ZN(n_0_194));
   NOR4_X1 i_0_244 (.A1(n_0_217), .A2(n_0_196), .A3(n_0_218), .A4(n_0_197), 
      .ZN(n_0_195));
   NAND4_X1 i_0_245 (.A1(n_0_338), .A2(n_0_346), .A3(n_0_332), .A4(n_0_341), 
      .ZN(n_0_196));
   AOI211_X1 i_0_246 (.A(n_0_203), .B(n_0_198), .C1(n_0_222), .C2(n_0_207), 
      .ZN(n_0_197));
   AOI21_X1 i_0_247 (.A(n_0_212), .B1(n_0_200), .B2(n_0_199), .ZN(n_0_198));
   NAND3_X1 i_0_248 (.A1(n_0_214), .A2(n_0_210), .A3(n_0_368), .ZN(n_0_199));
   NOR2_X1 i_0_249 (.A1(n_0_370), .A2(n_0_44), .ZN(n_0_200));
   NAND4_X1 i_0_250 (.A1(n_0_221), .A2(n_0_206), .A3(n_0_205), .A4(n_0_204), 
      .ZN(n_0_203));
   NAND2_X1 i_0_251 (.A1(i_add2[9]), .A2(i_add1[9]), .ZN(n_0_204));
   NAND2_X1 i_0_252 (.A1(i_add2[11]), .A2(i_add1[11]), .ZN(n_0_205));
   NAND2_X1 i_0_253 (.A1(i_add2[10]), .A2(i_add1[10]), .ZN(n_0_206));
   AND4_X1 i_0_254 (.A1(n_0_214), .A2(n_0_211), .A3(n_0_210), .A4(n_0_208), 
      .ZN(n_0_207));
   OR2_X1 i_0_255 (.A1(i_add2[5]), .A2(i_add1[5]), .ZN(n_0_208));
   OR2_X1 i_0_256 (.A1(i_add2[7]), .A2(i_add1[7]), .ZN(n_0_210));
   INV_X1 i_0_257 (.A(n_0_212), .ZN(n_0_211));
   NOR2_X1 i_0_258 (.A1(i_add2[8]), .A2(i_add1[8]), .ZN(n_0_212));
   OR2_X1 i_0_259 (.A1(i_add2[6]), .A2(i_add1[6]), .ZN(n_0_214));
   INV_X1 i_0_260 (.A(n_0_217), .ZN(n_0_215));
   NOR2_X1 i_0_261 (.A1(i_add2[13]), .A2(i_add1[13]), .ZN(n_0_217));
   INV_X1 i_0_262 (.A(n_0_220), .ZN(n_0_218));
   NAND3_X1 i_0_263 (.A1(n_0_360), .A2(n_0_221), .A3(n_0_361), .ZN(n_0_220));
   NAND2_X1 i_0_264 (.A1(i_add2[12]), .A2(i_add1[12]), .ZN(n_0_221));
   OAI21_X1 i_0_265 (.A(n_0_224), .B1(n_0_234), .B2(n_0_225), .ZN(n_0_222));
   NAND2_X1 i_0_266 (.A1(i_add2[5]), .A2(i_add1[5]), .ZN(n_0_224));
   AOI21_X1 i_0_267 (.A(n_0_373), .B1(n_0_375), .B2(n_0_374), .ZN(n_0_225));
   NOR2_X1 i_0_268 (.A1(i_add2[52]), .A2(i_add1[52]), .ZN(n_0_226));
   INV_X1 i_0_269 (.A(n_0_38), .ZN(n_0_227));
   INV_X1 i_0_270 (.A(n_0_39), .ZN(n_0_228));
   INV_X1 i_0_271 (.A(n_0_50), .ZN(n_0_229));
   INV_X1 i_0_272 (.A(n_0_42), .ZN(n_0_234));
   INV_X1 i_0_273 (.A(i_add1[43]), .ZN(n_0_236));
   INV_X1 i_0_274 (.A(i_add2[43]), .ZN(n_0_239));
   AOI21_X1 i_0_275 (.A(n_0_250), .B1(n_0_148), .B2(n_0_241), .ZN(n_0_240));
   OAI22_X1 i_0_276 (.A1(i_add2[37]), .A2(i_add1[37]), .B1(n_0_248), .B2(n_0_242), 
      .ZN(n_0_241));
   NAND2_X1 i_0_277 (.A1(n_0_164), .A2(n_0_243), .ZN(n_0_242));
   NAND3_X1 i_0_278 (.A1(n_0_102), .A2(n_0_244), .A3(n_0_108), .ZN(n_0_243));
   NAND2_X1 i_0_279 (.A1(n_0_150), .A2(n_0_245), .ZN(n_0_244));
   AOI21_X1 i_0_280 (.A(n_0_160), .B1(n_0_249), .B2(n_0_246), .ZN(n_0_245));
   NOR2_X1 i_0_281 (.A1(n_0_134), .A2(n_0_247), .ZN(n_0_246));
   NOR2_X1 i_0_282 (.A1(n_0_195), .A2(n_0_165), .ZN(n_0_247));
   INV_X1 i_0_283 (.A(n_0_149), .ZN(n_0_248));
   INV_X1 i_0_284 (.A(n_0_118), .ZN(n_0_249));
   INV_X1 i_0_285 (.A(n_0_89), .ZN(n_0_250));
   AOI21_X1 i_0_286 (.A(n_0_260), .B1(n_0_175), .B2(n_0_252), .ZN(n_0_251));
   NAND2_X1 i_0_287 (.A1(n_0_255), .A2(n_0_253), .ZN(n_0_252));
   OAI21_X1 i_0_288 (.A(n_0_177), .B1(n_0_257), .B2(n_0_254), .ZN(n_0_253));
   NOR3_X1 i_0_289 (.A1(n_0_265), .A2(n_0_195), .A3(n_0_184), .ZN(n_0_254));
   OR2_X1 i_0_290 (.A1(i_add2[17]), .A2(i_add1[17]), .ZN(n_0_255));
   INV_X1 i_0_291 (.A(n_0_257), .ZN(n_0_256));
   NOR2_X1 i_0_292 (.A1(i_add2[16]), .A2(i_add1[16]), .ZN(n_0_257));
   INV_X1 i_0_293 (.A(n_0_260), .ZN(n_0_258));
   NOR2_X1 i_0_294 (.A1(i_add2[18]), .A2(i_add1[18]), .ZN(n_0_260));
   INV_X1 i_0_295 (.A(n_0_179), .ZN(n_0_265));
   NAND2_X1 i_0_296 (.A1(n_0_269), .A2(n_0_266), .ZN(n_46));
   OAI221_X1 i_0_297 (.A(n_0_270), .B1(i_add2[62]), .B2(i_add1[62]), .C1(n_0_306), 
      .C2(n_0_267), .ZN(n_0_266));
   NOR2_X1 i_0_298 (.A1(n_0_271), .A2(n_0_268), .ZN(n_0_267));
   NOR3_X1 i_0_299 (.A1(n_0_282), .A2(n_0_279), .A3(n_0_275), .ZN(n_0_268));
   NAND2_X1 i_0_300 (.A1(i_add2[62]), .A2(i_add1[62]), .ZN(n_0_269));
   OR2_X1 i_0_301 (.A1(i_add2[61]), .A2(i_add1[61]), .ZN(n_0_270));
   OAI21_X1 i_0_302 (.A(n_0_272), .B1(i_add2[60]), .B2(i_add1[60]), .ZN(n_0_271));
   OAI21_X1 i_0_303 (.A(n_0_276), .B1(n_0_274), .B2(n_0_273), .ZN(n_0_272));
   NOR2_X1 i_0_304 (.A1(i_add2[58]), .A2(i_add1[58]), .ZN(n_0_273));
   NOR2_X1 i_0_305 (.A1(i_add2[59]), .A2(i_add1[59]), .ZN(n_0_274));
   OAI21_X1 i_0_306 (.A(n_0_276), .B1(n_0_314), .B2(n_0_311), .ZN(n_0_275));
   AOI21_X1 i_0_307 (.A(n_0_278), .B1(i_add2[60]), .B2(i_add1[60]), .ZN(n_0_276));
   NOR2_X1 i_0_308 (.A1(n_0_314), .A2(n_0_311), .ZN(n_0_277));
   AND2_X1 i_0_309 (.A1(i_add2[59]), .A2(i_add1[59]), .ZN(n_0_278));
   OAI22_X1 i_0_310 (.A1(n_0_313), .A2(n_0_310), .B1(n_0_288), .B2(n_0_280), 
      .ZN(n_0_279));
   AOI21_X1 i_0_311 (.A(n_0_281), .B1(i_add2[56]), .B2(i_add1[56]), .ZN(n_0_280));
   NOR2_X1 i_0_312 (.A1(n_0_312), .A2(n_0_309), .ZN(n_0_281));
   NOR3_X1 i_0_313 (.A1(n_0_287), .A2(n_0_283), .A3(n_0_296), .ZN(n_0_282));
   AOI22_X1 i_0_314 (.A1(i_add2[54]), .A2(i_add1[54]), .B1(n_0_286), .B2(n_0_284), 
      .ZN(n_0_283));
   OAI21_X1 i_0_315 (.A(n_0_305), .B1(n_0_226), .B2(n_0_285), .ZN(n_0_284));
   NOR3_X1 i_0_316 (.A1(i_add2[51]), .A2(n_0_308), .A3(i_add1[51]), .ZN(n_0_285));
   OR2_X1 i_0_317 (.A1(i_add2[53]), .A2(i_add1[53]), .ZN(n_0_286));
   NAND3_X1 i_0_318 (.A1(n_0_292), .A2(n_0_291), .A3(n_0_289), .ZN(n_0_287));
   INV_X1 i_0_319 (.A(n_0_289), .ZN(n_0_288));
   AOI21_X1 i_0_320 (.A(n_0_290), .B1(n_0_313), .B2(n_0_310), .ZN(n_0_289));
   NOR2_X1 i_0_321 (.A1(i_add2[56]), .A2(i_add1[56]), .ZN(n_0_290));
   NAND2_X1 i_0_322 (.A1(n_0_312), .A2(n_0_309), .ZN(n_0_291));
   OR2_X1 i_0_323 (.A1(i_add2[54]), .A2(i_add1[54]), .ZN(n_0_292));
   INV_X1 i_0_324 (.A(n_0_297), .ZN(n_0_296));
   NAND3_X1 i_0_325 (.A1(n_0_68), .A2(n_0_302), .A3(n_0_59), .ZN(n_0_297));
   INV_X1 i_0_326 (.A(n_0_303), .ZN(n_0_302));
   NAND3_X1 i_0_327 (.A1(n_0_56), .A2(n_0_305), .A3(n_0_304), .ZN(n_0_303));
   AOI21_X1 i_0_328 (.A(n_0_308), .B1(i_add2[54]), .B2(i_add1[54]), .ZN(n_0_304));
   NAND2_X1 i_0_329 (.A1(i_add2[53]), .A2(i_add1[53]), .ZN(n_0_305));
   INV_X1 i_0_330 (.A(n_0_307), .ZN(n_0_306));
   NAND2_X1 i_0_331 (.A1(i_add2[61]), .A2(i_add1[61]), .ZN(n_0_307));
   INV_X1 i_0_332 (.A(n_0_53), .ZN(n_0_308));
   INV_X1 i_0_333 (.A(i_add1[55]), .ZN(n_0_309));
   INV_X1 i_0_334 (.A(i_add1[57]), .ZN(n_0_310));
   INV_X1 i_0_335 (.A(i_add1[58]), .ZN(n_0_311));
   INV_X1 i_0_336 (.A(i_add2[55]), .ZN(n_0_312));
   INV_X1 i_0_337 (.A(i_add2[57]), .ZN(n_0_313));
   INV_X1 i_0_338 (.A(i_add2[58]), .ZN(n_0_314));
   OR2_X1 i_0_339 (.A1(n_0_283), .A2(n_0_287), .ZN(n_0_315));
   NOR2_X1 i_0_340 (.A1(n_0_279), .A2(n_0_275), .ZN(n_0_316));
   AND3_X1 i_0_341 (.A1(n_0_99), .A2(n_0_69), .A3(n_0_124), .ZN(n_0_317));
   NOR3_X1 i_0_342 (.A1(n_0_317), .A2(n_0_58), .A3(n_0_303), .ZN(n_0_318));
   AOI221_X1 i_0_343 (.A(n_0_271), .B1(n_0_315), .B2(n_0_316), .C1(n_0_318), 
      .C2(n_0_316), .ZN(n_0_319));
   INV_X1 i_0_344 (.A(n_0_270), .ZN(n_0_320));
   INV_X1 i_0_345 (.A(n_0_319), .ZN(n_0_321));
   AOI21_X1 i_0_346 (.A(n_0_320), .B1(n_0_321), .B2(n_0_307), .ZN(n_47));
   NOR2_X1 i_0_347 (.A1(n_0_274), .A2(n_0_322), .ZN(n_48));
   NOR2_X1 i_0_348 (.A1(n_0_278), .A2(n_0_323), .ZN(n_0_322));
   NOR2_X1 i_0_349 (.A1(n_0_273), .A2(n_0_324), .ZN(n_0_323));
   NOR3_X1 i_0_350 (.A1(n_0_279), .A2(n_0_277), .A3(n_0_282), .ZN(n_0_324));
   OR2_X1 i_0_351 (.A1(n_0_282), .A2(n_0_279), .ZN(n_49));
   NOR2_X1 i_0_352 (.A1(n_0_88), .A2(n_0_325), .ZN(n_50));
   NOR2_X1 i_0_353 (.A1(n_0_240), .A2(n_0_129), .ZN(n_0_325));
   INV_X1 i_0_354 (.A(n_51), .ZN(n_0_326));
   AOI21_X1 i_0_355 (.A(n_0_105), .B1(n_0_159), .B2(n_0_327), .ZN(n_51));
   INV_X1 i_0_356 (.A(n_0_328), .ZN(n_0_327));
   AOI21_X1 i_0_357 (.A(n_0_228), .B1(n_0_245), .B2(n_0_158), .ZN(n_0_328));
   AOI21_X1 i_0_358 (.A(n_0_257), .B1(n_0_179), .B2(n_0_329), .ZN(n_52));
   OAI21_X1 i_0_359 (.A(n_0_346), .B1(n_0_344), .B2(n_0_330), .ZN(n_0_329));
   NAND2_X1 i_0_360 (.A1(n_0_187), .A2(n_0_331), .ZN(n_0_330));
   NAND3_X1 i_0_361 (.A1(n_0_215), .A2(n_0_332), .A3(n_0_334), .ZN(n_0_331));
   INV_X1 i_0_362 (.A(n_0_333), .ZN(n_0_332));
   NOR2_X1 i_0_363 (.A1(i_add2[14]), .A2(i_add1[14]), .ZN(n_0_333));
   OAI21_X1 i_0_364 (.A(n_0_336), .B1(n_0_337), .B2(n_0_335), .ZN(n_0_334));
   OAI211_X1 i_0_365 (.A(n_0_220), .B(n_0_341), .C1(n_0_203), .C2(n_0_342), 
      .ZN(n_0_335));
   NAND2_X1 i_0_366 (.A1(i_add2[13]), .A2(i_add1[13]), .ZN(n_0_336));
   INV_X1 i_0_367 (.A(n_0_338), .ZN(n_0_337));
   OAI211_X1 i_0_368 (.A(n_0_205), .B(n_0_221), .C1(n_0_340), .C2(n_0_339), 
      .ZN(n_0_338));
   NOR3_X1 i_0_369 (.A1(i_add2[9]), .A2(n_0_347), .A3(i_add1[9]), .ZN(n_0_339));
   NOR2_X1 i_0_370 (.A1(i_add2[10]), .A2(i_add1[10]), .ZN(n_0_340));
   OR2_X1 i_0_371 (.A1(i_add2[12]), .A2(i_add1[12]), .ZN(n_0_341));
   INV_X1 i_0_372 (.A(n_0_343), .ZN(n_0_342));
   AOI21_X1 i_0_373 (.A(n_0_198), .B1(n_0_222), .B2(n_0_207), .ZN(n_0_343));
   INV_X1 i_0_374 (.A(n_0_345), .ZN(n_0_344));
   NAND2_X1 i_0_375 (.A1(i_add2[14]), .A2(i_add1[14]), .ZN(n_0_345));
   INV_X1 i_0_376 (.A(n_0_188), .ZN(n_0_346));
   INV_X1 i_0_377 (.A(n_0_206), .ZN(n_0_347));
   AND2_X1 i_0_378 (.A1(n_0_346), .A2(n_0_348), .ZN(n_53));
   OAI21_X1 i_0_379 (.A(n_0_187), .B1(n_0_333), .B2(n_0_349), .ZN(n_0_348));
   AOI21_X1 i_0_380 (.A(n_0_350), .B1(n_0_334), .B2(n_0_215), .ZN(n_0_349));
   INV_X1 i_0_381 (.A(n_0_345), .ZN(n_0_350));
   AND2_X1 i_0_382 (.A1(n_0_215), .A2(n_0_351), .ZN(n_54));
   OAI21_X1 i_0_383 (.A(n_0_336), .B1(n_0_358), .B2(n_0_352), .ZN(n_0_351));
   AOI21_X1 i_0_384 (.A(n_0_359), .B1(n_0_355), .B2(n_0_353), .ZN(n_0_352));
   OAI21_X1 i_0_385 (.A(n_0_205), .B1(n_0_340), .B2(n_0_354), .ZN(n_0_353));
   AOI21_X1 i_0_386 (.A(n_0_347), .B1(n_0_357), .B2(n_0_356), .ZN(n_0_354));
   NAND2_X1 i_0_387 (.A1(n_0_361), .A2(n_0_360), .ZN(n_0_355));
   OR2_X1 i_0_388 (.A1(i_add1[9]), .A2(i_add2[9]), .ZN(n_0_356));
   NAND2_X1 i_0_389 (.A1(n_0_343), .A2(n_0_204), .ZN(n_0_357));
   INV_X1 i_0_390 (.A(n_0_341), .ZN(n_0_358));
   INV_X1 i_0_391 (.A(n_0_221), .ZN(n_0_359));
   INV_X1 i_0_392 (.A(i_add2[11]), .ZN(n_0_360));
   INV_X1 i_0_393 (.A(i_add1[11]), .ZN(n_0_361));
   AND2_X1 i_0_394 (.A1(n_0_355), .A2(n_0_362), .ZN(n_55));
   OAI21_X1 i_0_395 (.A(n_0_205), .B1(n_0_340), .B2(n_0_363), .ZN(n_0_362));
   AOI21_X1 i_0_396 (.A(n_0_364), .B1(n_0_356), .B2(n_0_43), .ZN(n_0_363));
   INV_X1 i_0_397 (.A(n_0_206), .ZN(n_0_364));
   AND2_X1 i_0_398 (.A1(n_0_43), .A2(n_0_356), .ZN(n_56));
   NOR2_X1 i_0_399 (.A1(n_0_371), .A2(n_0_365), .ZN(n_57));
   AOI21_X1 i_0_400 (.A(n_0_370), .B1(n_0_210), .B2(n_0_366), .ZN(n_0_365));
   OAI21_X1 i_0_401 (.A(n_0_369), .B1(n_0_372), .B2(n_0_367), .ZN(n_0_366));
   AOI21_X1 i_0_402 (.A(n_0_368), .B1(n_0_222), .B2(n_0_208), .ZN(n_0_367));
   AND2_X1 i_0_403 (.A1(i_add1[6]), .A2(i_add2[6]), .ZN(n_0_368));
   NAND2_X1 i_0_404 (.A1(i_add1[7]), .A2(i_add2[7]), .ZN(n_0_369));
   AND2_X1 i_0_405 (.A1(i_add1[8]), .A2(i_add2[8]), .ZN(n_0_370));
   INV_X1 i_0_406 (.A(n_0_211), .ZN(n_0_371));
   INV_X1 i_0_407 (.A(n_0_214), .ZN(n_0_372));
   AND2_X1 i_0_408 (.A1(n_0_366), .A2(n_0_210), .ZN(n_58));
   AND2_X1 i_0_409 (.A1(n_0_222), .A2(n_0_208), .ZN(n_59));
   AND2_X1 i_0_410 (.A1(i_add2[4]), .A2(i_add1[4]), .ZN(n_0_373));
   AND2_X1 i_0_411 (.A1(n_0_375), .A2(n_0_374), .ZN(n_60));
   NAND2_X1 i_0_412 (.A1(n_0_383), .A2(n_0_382), .ZN(n_0_374));
   OAI22_X1 i_0_413 (.A1(n_0_383), .A2(n_0_382), .B1(n_0_377), .B2(n_0_376), 
      .ZN(n_0_375));
   NOR2_X1 i_0_414 (.A1(i_add2[2]), .A2(i_add1[2]), .ZN(n_0_376));
   AOI22_X1 i_0_415 (.A1(n_0_379), .A2(n_0_378), .B1(i_add2[2]), .B2(i_add1[2]), 
      .ZN(n_0_377));
   OR2_X1 i_0_416 (.A1(i_add2[1]), .A2(i_add1[1]), .ZN(n_0_378));
   NAND2_X1 i_0_417 (.A1(n_0_381), .A2(n_0_380), .ZN(n_0_379));
   NAND2_X1 i_0_418 (.A1(i_add2[1]), .A2(i_add1[1]), .ZN(n_0_380));
   NAND2_X1 i_0_419 (.A1(i_add2[0]), .A2(i_add1[0]), .ZN(n_0_381));
   INV_X1 i_0_420 (.A(i_add1[3]), .ZN(n_0_382));
   INV_X1 i_0_421 (.A(i_add2[3]), .ZN(n_0_383));
   AND2_X1 i_0_422 (.A1(n_0_379), .A2(n_0_378), .ZN(n_61));
endmodule

module regFile64(read_data, write_en, write_data, clk);
   output [63:0]read_data;
   input write_en;
   input [63:0]write_data;
   input clk;

   DFF_X1 \my_reg_reg[63]  (.D(write_data[63]), .CK(n_0), .Q(read_data[63]), 
      .QN());
   INV_X1 i_0_0 (.A(clk), .ZN(n_0));
   DFF_X1 \my_reg_reg[62]  (.D(write_data[62]), .CK(n_0), .Q(read_data[62]), 
      .QN());
   DFF_X1 \my_reg_reg[61]  (.D(write_data[61]), .CK(n_0), .Q(read_data[61]), 
      .QN());
   DFF_X1 \my_reg_reg[60]  (.D(write_data[60]), .CK(n_0), .Q(read_data[60]), 
      .QN());
   DFF_X1 \my_reg_reg[59]  (.D(write_data[59]), .CK(n_0), .Q(read_data[59]), 
      .QN());
   DFF_X1 \my_reg_reg[58]  (.D(write_data[58]), .CK(n_0), .Q(read_data[58]), 
      .QN());
   DFF_X1 \my_reg_reg[57]  (.D(write_data[57]), .CK(n_0), .Q(read_data[57]), 
      .QN());
   DFF_X1 \my_reg_reg[56]  (.D(write_data[56]), .CK(n_0), .Q(read_data[56]), 
      .QN());
   DFF_X1 \my_reg_reg[55]  (.D(write_data[55]), .CK(n_0), .Q(read_data[55]), 
      .QN());
   DFF_X1 \my_reg_reg[54]  (.D(write_data[54]), .CK(n_0), .Q(read_data[54]), 
      .QN());
   DFF_X1 \my_reg_reg[53]  (.D(write_data[53]), .CK(n_0), .Q(read_data[53]), 
      .QN());
   DFF_X1 \my_reg_reg[52]  (.D(write_data[52]), .CK(n_0), .Q(read_data[52]), 
      .QN());
   DFF_X1 \my_reg_reg[51]  (.D(write_data[51]), .CK(n_0), .Q(read_data[51]), 
      .QN());
   DFF_X1 \my_reg_reg[50]  (.D(write_data[50]), .CK(n_0), .Q(read_data[50]), 
      .QN());
   DFF_X1 \my_reg_reg[49]  (.D(write_data[49]), .CK(n_0), .Q(read_data[49]), 
      .QN());
   DFF_X1 \my_reg_reg[48]  (.D(write_data[48]), .CK(n_0), .Q(read_data[48]), 
      .QN());
   DFF_X1 \my_reg_reg[47]  (.D(write_data[47]), .CK(n_0), .Q(read_data[47]), 
      .QN());
   DFF_X1 \my_reg_reg[46]  (.D(write_data[46]), .CK(n_0), .Q(read_data[46]), 
      .QN());
   DFF_X1 \my_reg_reg[45]  (.D(write_data[45]), .CK(n_0), .Q(read_data[45]), 
      .QN());
   DFF_X1 \my_reg_reg[44]  (.D(write_data[44]), .CK(n_0), .Q(read_data[44]), 
      .QN());
   DFF_X1 \my_reg_reg[43]  (.D(write_data[43]), .CK(n_0), .Q(read_data[43]), 
      .QN());
   DFF_X1 \my_reg_reg[42]  (.D(write_data[42]), .CK(n_0), .Q(read_data[42]), 
      .QN());
   DFF_X1 \my_reg_reg[41]  (.D(write_data[41]), .CK(n_0), .Q(read_data[41]), 
      .QN());
   DFF_X1 \my_reg_reg[40]  (.D(write_data[40]), .CK(n_0), .Q(read_data[40]), 
      .QN());
   DFF_X1 \my_reg_reg[39]  (.D(write_data[39]), .CK(n_0), .Q(read_data[39]), 
      .QN());
   DFF_X1 \my_reg_reg[38]  (.D(write_data[38]), .CK(n_0), .Q(read_data[38]), 
      .QN());
   DFF_X1 \my_reg_reg[37]  (.D(write_data[37]), .CK(n_0), .Q(read_data[37]), 
      .QN());
   DFF_X1 \my_reg_reg[36]  (.D(write_data[36]), .CK(n_0), .Q(read_data[36]), 
      .QN());
   DFF_X1 \my_reg_reg[35]  (.D(write_data[35]), .CK(n_0), .Q(read_data[35]), 
      .QN());
   DFF_X1 \my_reg_reg[34]  (.D(write_data[34]), .CK(n_0), .Q(read_data[34]), 
      .QN());
   DFF_X1 \my_reg_reg[33]  (.D(write_data[33]), .CK(n_0), .Q(read_data[33]), 
      .QN());
   DFF_X1 \my_reg_reg[32]  (.D(write_data[32]), .CK(n_0), .Q(read_data[32]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
endmodule

module datapath__0_193(p_0, read_data2);
   output [31:0]p_0;
   input [31:0]read_data2;

   XOR2_X1 i_0 (.A(read_data2[1]), .B(read_data2[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(read_data2[2]), .B1(read_data2[1]), .B2(read_data2[0]), 
      .ZN(n_0));
   XOR2_X1 i_3 (.A(read_data2[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(read_data2[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(read_data2[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(read_data2[6]), .B1(n_27), .B2(read_data2[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(read_data2[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(read_data2[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(read_data2[9]), .B1(n_25), .B2(read_data2[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(read_data2[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(read_data2[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(read_data2[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(read_data2[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(read_data2[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(read_data2[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(read_data2[16]), .B1(n_19), .B2(read_data2[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(read_data2[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(read_data2[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(read_data2[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(read_data2[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(read_data2[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(read_data2[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(read_data2[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(read_data2[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(read_data2[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(read_data2[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(read_data2[27]), .B1(n_9), .B2(read_data2[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(read_data2[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(read_data2[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(read_data2[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(read_data2[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(read_data2[28]), .A3(read_data2[29]), .A4(
      read_data2[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(read_data2[28]), .A3(read_data2[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(read_data2[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(read_data2[26]), .A3(read_data2[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(read_data2[23]), .A3(read_data2[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(read_data2[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(read_data2[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(read_data2[18]), .A3(read_data2[19]), .A4(
      read_data2[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(read_data2[18]), .A3(read_data2[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(read_data2[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(read_data2[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(read_data2[15]), .A3(read_data2[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(read_data2[12]), .A3(read_data2[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(read_data2[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(read_data2[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(read_data2[8]), .A3(read_data2[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(read_data2[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(read_data2[5]), .A3(read_data2[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(read_data2[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(read_data2[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(read_data2[2]), .A2(read_data2[1]), .A3(read_data2[0]), 
      .ZN(n_29));
   INV_X1 i_61 (.A(read_data2[11]), .ZN(n_30));
   INV_X1 i_62 (.A(read_data2[14]), .ZN(n_31));
   INV_X1 i_63 (.A(read_data2[21]), .ZN(n_32));
   INV_X1 i_64 (.A(read_data2[25]), .ZN(n_33));
endmodule

module datapath__0_195(p_0, p_1);
   output [32:0]p_0;
   input [32:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_27), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_25), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(p_1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(p_1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(p_1[16]), .B1(n_19), .B2(p_1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(p_1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(p_1[27]), .B1(n_9), .B2(p_1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(p_1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(p_1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(p_1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(p_1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(p_1[26]), .A3(p_1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(p_1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(p_1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(p_1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(p_1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(p_1[15]), .A3(p_1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(p_1[12]), .A3(p_1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(p_1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(p_1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(p_1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(p_1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(p_1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(p_1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(p_1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(p_1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(p_1[25]), .ZN(n_33));
endmodule

module Radix4(a, b, read_data3, clk, start, start_shift, start_i);
   input [31:0]a;
   input [31:0]b;
   output [63:0]read_data3;
   input clk;
   input start;
   input [4:0]start_shift;
   input [4:0]start_i;

   wire [31:0]read_data2;
   wire [31:0]read_data;
   wire [63:0]res;
   wire [63:0]sum;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_0_0;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_0_1;
   wire n_0_126;
   wire n_0_0_2;
   wire n_0_127;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_128;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_129;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_130;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_131;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_176;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_177;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_178;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_179;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_180;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_181;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_182;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_183;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_184;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_185;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_186;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_187;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_188;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_189;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_190;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_191;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_192;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_193;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_194;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_195;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_196;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_197;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_198;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_199;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_200;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_201;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_132;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_133;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_134;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_135;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_136;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_137;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_138;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_139;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_140;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_141;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_142;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_143;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_144;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_145;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_146;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_147;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_148;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_149;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_150;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_151;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_152;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_153;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_154;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_155;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_156;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_157;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_158;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_159;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_160;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_161;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_162;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_163;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_164;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_165;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_166;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_167;
   wire n_0_169;
   wire n_0_0_442;
   wire n_0_168;
   wire n_0_0_443;
   wire n_0_170;
   wire n_0_0_444;
   wire n_0_171;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_172;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_173;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_174;
   wire write_en;
   wire [63:0]c;
   wire [4:0]shift;
   wire [4:0]i;
   wire n_0_175;

   regFile r (.read_data(read_data), .read_data2(read_data2), .write_en(write_en), 
      .write_data(a), .write_data2(b), .clk(clk));
   carry_lookahead_adder ADD (.i_add1(c), .i_add2(sum), .o_result(res), .o_carry());
   regFile64 r2 (.read_data(read_data3), .write_en(), .write_data(res), .clk(clk));
   DFF_X1 \sum_reg[63]  (.D(n_0_169), .CK(clk), .Q(sum[63]), .QN());
   DFF_X1 \sum_reg[62]  (.D(n_0_168), .CK(clk), .Q(sum[62]), .QN());
   DFF_X1 \sum_reg[61]  (.D(n_0_167), .CK(clk), .Q(sum[61]), .QN());
   DFF_X1 \sum_reg[60]  (.D(n_0_166), .CK(clk), .Q(sum[60]), .QN());
   DFF_X1 \sum_reg[59]  (.D(n_0_165), .CK(clk), .Q(sum[59]), .QN());
   DFF_X1 \sum_reg[58]  (.D(n_0_164), .CK(clk), .Q(sum[58]), .QN());
   DFF_X1 \sum_reg[57]  (.D(n_0_163), .CK(clk), .Q(sum[57]), .QN());
   DFF_X1 \sum_reg[56]  (.D(n_0_162), .CK(clk), .Q(sum[56]), .QN());
   DFF_X1 \sum_reg[55]  (.D(n_0_161), .CK(clk), .Q(sum[55]), .QN());
   DFF_X1 \sum_reg[54]  (.D(n_0_160), .CK(clk), .Q(sum[54]), .QN());
   DFF_X1 \sum_reg[53]  (.D(n_0_159), .CK(clk), .Q(sum[53]), .QN());
   DFF_X1 \sum_reg[52]  (.D(n_0_158), .CK(clk), .Q(sum[52]), .QN());
   DFF_X1 \sum_reg[51]  (.D(n_0_157), .CK(clk), .Q(sum[51]), .QN());
   DFF_X1 \sum_reg[50]  (.D(n_0_156), .CK(clk), .Q(sum[50]), .QN());
   DFF_X1 \sum_reg[49]  (.D(n_0_155), .CK(clk), .Q(sum[49]), .QN());
   DFF_X1 \sum_reg[48]  (.D(n_0_154), .CK(clk), .Q(sum[48]), .QN());
   DFF_X1 \sum_reg[47]  (.D(n_0_153), .CK(clk), .Q(sum[47]), .QN());
   DFF_X1 \sum_reg[46]  (.D(n_0_152), .CK(clk), .Q(sum[46]), .QN());
   DFF_X1 \sum_reg[45]  (.D(n_0_151), .CK(clk), .Q(sum[45]), .QN());
   DFF_X1 \sum_reg[44]  (.D(n_0_150), .CK(clk), .Q(sum[44]), .QN());
   DFF_X1 \sum_reg[43]  (.D(n_0_149), .CK(clk), .Q(sum[43]), .QN());
   DFF_X1 \sum_reg[42]  (.D(n_0_148), .CK(clk), .Q(sum[42]), .QN());
   DFF_X1 \sum_reg[41]  (.D(n_0_147), .CK(clk), .Q(sum[41]), .QN());
   DFF_X1 \sum_reg[40]  (.D(n_0_146), .CK(clk), .Q(sum[40]), .QN());
   DFF_X1 \sum_reg[39]  (.D(n_0_145), .CK(clk), .Q(sum[39]), .QN());
   DFF_X1 \sum_reg[38]  (.D(n_0_144), .CK(clk), .Q(sum[38]), .QN());
   DFF_X1 \sum_reg[37]  (.D(n_0_143), .CK(clk), .Q(sum[37]), .QN());
   DFF_X1 \sum_reg[36]  (.D(n_0_142), .CK(clk), .Q(sum[36]), .QN());
   DFF_X1 \sum_reg[35]  (.D(n_0_141), .CK(clk), .Q(sum[35]), .QN());
   DFF_X1 \sum_reg[34]  (.D(n_0_140), .CK(clk), .Q(sum[34]), .QN());
   DFF_X1 \sum_reg[33]  (.D(n_0_139), .CK(clk), .Q(sum[33]), .QN());
   DFF_X1 \sum_reg[32]  (.D(n_0_138), .CK(clk), .Q(sum[32]), .QN());
   DFF_X1 \sum_reg[31]  (.D(n_0_137), .CK(clk), .Q(sum[31]), .QN());
   DFF_X1 \sum_reg[30]  (.D(n_0_136), .CK(clk), .Q(sum[30]), .QN());
   DFF_X1 \sum_reg[29]  (.D(n_0_135), .CK(clk), .Q(sum[29]), .QN());
   DFF_X1 \sum_reg[28]  (.D(n_0_134), .CK(clk), .Q(sum[28]), .QN());
   DFF_X1 \sum_reg[27]  (.D(n_0_133), .CK(clk), .Q(sum[27]), .QN());
   DFF_X1 \sum_reg[26]  (.D(n_0_132), .CK(clk), .Q(sum[26]), .QN());
   DFF_X1 \sum_reg[25]  (.D(n_0_201), .CK(clk), .Q(sum[25]), .QN());
   DFF_X1 \sum_reg[24]  (.D(n_0_200), .CK(clk), .Q(sum[24]), .QN());
   DFF_X1 \sum_reg[23]  (.D(n_0_199), .CK(clk), .Q(sum[23]), .QN());
   DFF_X1 \sum_reg[22]  (.D(n_0_198), .CK(clk), .Q(sum[22]), .QN());
   DFF_X1 \sum_reg[21]  (.D(n_0_197), .CK(clk), .Q(sum[21]), .QN());
   DFF_X1 \sum_reg[20]  (.D(n_0_196), .CK(clk), .Q(sum[20]), .QN());
   DFF_X1 \sum_reg[19]  (.D(n_0_195), .CK(clk), .Q(sum[19]), .QN());
   DFF_X1 \sum_reg[18]  (.D(n_0_194), .CK(clk), .Q(sum[18]), .QN());
   DFF_X1 \sum_reg[17]  (.D(n_0_193), .CK(clk), .Q(sum[17]), .QN());
   DFF_X1 \sum_reg[16]  (.D(n_0_192), .CK(clk), .Q(sum[16]), .QN());
   DFF_X1 \sum_reg[15]  (.D(n_0_191), .CK(clk), .Q(sum[15]), .QN());
   DFF_X1 \sum_reg[14]  (.D(n_0_190), .CK(clk), .Q(sum[14]), .QN());
   DFF_X1 \sum_reg[13]  (.D(n_0_189), .CK(clk), .Q(sum[13]), .QN());
   DFF_X1 \sum_reg[12]  (.D(n_0_188), .CK(clk), .Q(sum[12]), .QN());
   DFF_X1 \sum_reg[11]  (.D(n_0_187), .CK(clk), .Q(sum[11]), .QN());
   DFF_X1 \sum_reg[10]  (.D(n_0_186), .CK(clk), .Q(sum[10]), .QN());
   DFF_X1 \sum_reg[9]  (.D(n_0_185), .CK(clk), .Q(sum[9]), .QN());
   DFF_X1 \sum_reg[8]  (.D(n_0_184), .CK(clk), .Q(sum[8]), .QN());
   DFF_X1 \sum_reg[7]  (.D(n_0_183), .CK(clk), .Q(sum[7]), .QN());
   DFF_X1 \sum_reg[6]  (.D(n_0_182), .CK(clk), .Q(sum[6]), .QN());
   DFF_X1 \sum_reg[5]  (.D(n_0_181), .CK(clk), .Q(sum[5]), .QN());
   DFF_X1 \sum_reg[4]  (.D(n_0_180), .CK(clk), .Q(sum[4]), .QN());
   DFF_X1 \sum_reg[3]  (.D(n_0_179), .CK(clk), .Q(sum[3]), .QN());
   DFF_X1 \sum_reg[2]  (.D(n_0_178), .CK(clk), .Q(sum[2]), .QN());
   DFF_X1 \sum_reg[1]  (.D(n_0_177), .CK(clk), .Q(sum[1]), .QN());
   DFF_X1 \sum_reg[0]  (.D(n_0_176), .CK(clk), .Q(sum[0]), .QN());
   datapath__0_193 i_0_2 (.p_0({n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, 
      n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, uc_0}), .read_data2(
      read_data2));
   datapath__0_195 i_0_3 (.p_0({uc_1, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, 
      n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, 
      n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, uc_2}), 
      .p_1({1'b0, read_data2[31], read_data2[30], read_data2[29], read_data2[28], 
      read_data2[27], read_data2[26], read_data2[25], read_data2[24], 
      read_data2[23], read_data2[22], read_data2[21], read_data2[20], 
      read_data2[19], read_data2[18], read_data2[17], read_data2[16], 
      read_data2[15], read_data2[14], read_data2[13], read_data2[12], 
      read_data2[11], read_data2[10], read_data2[9], read_data2[8], 
      read_data2[7], read_data2[6], read_data2[5], read_data2[4], read_data2[3], 
      read_data2[2], read_data2[1], read_data2[0]}));
   INV_X1 i_0_0_0 (.A(start), .ZN(n_0_0_0));
   AND2_X1 i_0_0_1 (.A1(n_0_0_0), .A2(res[0]), .ZN(n_0_0));
   AND2_X1 i_0_0_2 (.A1(n_0_0_0), .A2(res[1]), .ZN(n_0_1));
   AND2_X1 i_0_0_3 (.A1(n_0_0_0), .A2(res[2]), .ZN(n_0_2));
   AND2_X1 i_0_0_4 (.A1(n_0_0_0), .A2(res[3]), .ZN(n_0_3));
   AND2_X1 i_0_0_5 (.A1(n_0_0_0), .A2(res[4]), .ZN(n_0_4));
   AND2_X1 i_0_0_6 (.A1(n_0_0_0), .A2(res[5]), .ZN(n_0_5));
   AND2_X1 i_0_0_7 (.A1(n_0_0_0), .A2(res[6]), .ZN(n_0_6));
   AND2_X1 i_0_0_8 (.A1(n_0_0_0), .A2(res[7]), .ZN(n_0_7));
   AND2_X1 i_0_0_9 (.A1(n_0_0_0), .A2(res[8]), .ZN(n_0_8));
   AND2_X1 i_0_0_10 (.A1(n_0_0_0), .A2(res[9]), .ZN(n_0_71));
   AND2_X1 i_0_0_11 (.A1(n_0_0_0), .A2(res[10]), .ZN(n_0_72));
   AND2_X1 i_0_0_12 (.A1(n_0_0_0), .A2(res[11]), .ZN(n_0_73));
   AND2_X1 i_0_0_13 (.A1(n_0_0_0), .A2(res[12]), .ZN(n_0_74));
   AND2_X1 i_0_0_14 (.A1(n_0_0_0), .A2(res[13]), .ZN(n_0_75));
   AND2_X1 i_0_0_15 (.A1(n_0_0_0), .A2(res[14]), .ZN(n_0_76));
   AND2_X1 i_0_0_16 (.A1(n_0_0_0), .A2(res[15]), .ZN(n_0_77));
   AND2_X1 i_0_0_17 (.A1(n_0_0_0), .A2(res[16]), .ZN(n_0_78));
   AND2_X1 i_0_0_18 (.A1(n_0_0_0), .A2(res[17]), .ZN(n_0_79));
   AND2_X1 i_0_0_19 (.A1(n_0_0_0), .A2(res[18]), .ZN(n_0_80));
   AND2_X1 i_0_0_20 (.A1(n_0_0_0), .A2(res[19]), .ZN(n_0_81));
   AND2_X1 i_0_0_21 (.A1(n_0_0_0), .A2(res[20]), .ZN(n_0_82));
   AND2_X1 i_0_0_22 (.A1(n_0_0_0), .A2(res[21]), .ZN(n_0_83));
   AND2_X1 i_0_0_23 (.A1(n_0_0_0), .A2(res[22]), .ZN(n_0_84));
   AND2_X1 i_0_0_24 (.A1(n_0_0_0), .A2(res[23]), .ZN(n_0_85));
   AND2_X1 i_0_0_25 (.A1(n_0_0_0), .A2(res[24]), .ZN(n_0_86));
   AND2_X1 i_0_0_26 (.A1(n_0_0_0), .A2(res[25]), .ZN(n_0_87));
   AND2_X1 i_0_0_27 (.A1(n_0_0_0), .A2(res[26]), .ZN(n_0_88));
   AND2_X1 i_0_0_28 (.A1(n_0_0_0), .A2(res[27]), .ZN(n_0_89));
   AND2_X1 i_0_0_29 (.A1(n_0_0_0), .A2(res[28]), .ZN(n_0_90));
   AND2_X1 i_0_0_30 (.A1(n_0_0_0), .A2(res[29]), .ZN(n_0_91));
   AND2_X1 i_0_0_31 (.A1(n_0_0_0), .A2(res[30]), .ZN(n_0_92));
   AND2_X1 i_0_0_32 (.A1(n_0_0_0), .A2(res[31]), .ZN(n_0_93));
   AND2_X1 i_0_0_33 (.A1(n_0_0_0), .A2(res[32]), .ZN(n_0_94));
   AND2_X1 i_0_0_34 (.A1(n_0_0_0), .A2(res[33]), .ZN(n_0_95));
   AND2_X1 i_0_0_35 (.A1(n_0_0_0), .A2(res[34]), .ZN(n_0_96));
   AND2_X1 i_0_0_36 (.A1(n_0_0_0), .A2(res[35]), .ZN(n_0_97));
   AND2_X1 i_0_0_37 (.A1(n_0_0_0), .A2(res[36]), .ZN(n_0_98));
   AND2_X1 i_0_0_38 (.A1(n_0_0_0), .A2(res[37]), .ZN(n_0_99));
   AND2_X1 i_0_0_39 (.A1(n_0_0_0), .A2(res[38]), .ZN(n_0_100));
   AND2_X1 i_0_0_40 (.A1(n_0_0_0), .A2(res[39]), .ZN(n_0_101));
   AND2_X1 i_0_0_41 (.A1(n_0_0_0), .A2(res[40]), .ZN(n_0_102));
   AND2_X1 i_0_0_42 (.A1(n_0_0_0), .A2(res[41]), .ZN(n_0_103));
   AND2_X1 i_0_0_43 (.A1(n_0_0_0), .A2(res[42]), .ZN(n_0_104));
   AND2_X1 i_0_0_44 (.A1(n_0_0_0), .A2(res[43]), .ZN(n_0_105));
   AND2_X1 i_0_0_45 (.A1(n_0_0_0), .A2(res[44]), .ZN(n_0_106));
   AND2_X1 i_0_0_46 (.A1(n_0_0_0), .A2(res[45]), .ZN(n_0_107));
   AND2_X1 i_0_0_47 (.A1(n_0_0_0), .A2(res[46]), .ZN(n_0_108));
   AND2_X1 i_0_0_48 (.A1(n_0_0_0), .A2(res[47]), .ZN(n_0_109));
   AND2_X1 i_0_0_49 (.A1(n_0_0_0), .A2(res[48]), .ZN(n_0_110));
   AND2_X1 i_0_0_50 (.A1(n_0_0_0), .A2(res[49]), .ZN(n_0_111));
   AND2_X1 i_0_0_51 (.A1(n_0_0_0), .A2(res[50]), .ZN(n_0_112));
   AND2_X1 i_0_0_52 (.A1(n_0_0_0), .A2(res[51]), .ZN(n_0_113));
   AND2_X1 i_0_0_53 (.A1(n_0_0_0), .A2(res[52]), .ZN(n_0_114));
   AND2_X1 i_0_0_54 (.A1(n_0_0_0), .A2(res[53]), .ZN(n_0_115));
   AND2_X1 i_0_0_55 (.A1(n_0_0_0), .A2(res[54]), .ZN(n_0_116));
   AND2_X1 i_0_0_56 (.A1(n_0_0_0), .A2(res[55]), .ZN(n_0_117));
   AND2_X1 i_0_0_57 (.A1(n_0_0_0), .A2(res[56]), .ZN(n_0_118));
   AND2_X1 i_0_0_58 (.A1(n_0_0_0), .A2(res[57]), .ZN(n_0_119));
   AND2_X1 i_0_0_59 (.A1(n_0_0_0), .A2(res[58]), .ZN(n_0_120));
   AND2_X1 i_0_0_60 (.A1(n_0_0_0), .A2(res[59]), .ZN(n_0_121));
   AND2_X1 i_0_0_61 (.A1(n_0_0_0), .A2(res[60]), .ZN(n_0_122));
   AND2_X1 i_0_0_62 (.A1(n_0_0_0), .A2(res[61]), .ZN(n_0_123));
   AND2_X1 i_0_0_63 (.A1(n_0_0_0), .A2(res[62]), .ZN(n_0_124));
   AND2_X1 i_0_0_64 (.A1(n_0_0_0), .A2(res[63]), .ZN(n_0_125));
   OAI22_X1 i_0_0_65 (.A1(n_0_0_0), .A2(start_i[0]), .B1(i[0]), .B2(start), 
      .ZN(n_0_0_1));
   INV_X1 i_0_0_66 (.A(n_0_0_1), .ZN(n_0_126));
   INV_X1 i_0_0_67 (.A(start_i[1]), .ZN(n_0_0_2));
   AOI22_X1 i_0_0_68 (.A1(n_0_0_2), .A2(start), .B1(n_0_0_0), .B2(i[1]), 
      .ZN(n_0_127));
   NAND2_X1 i_0_0_69 (.A1(start_i[2]), .A2(start), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_70 (.A(n_0_0_0), .B1(i[2]), .B2(i[1]), .ZN(n_0_0_4));
   NAND2_X1 i_0_0_71 (.A1(i[2]), .A2(i[1]), .ZN(n_0_0_5));
   INV_X1 i_0_0_72 (.A(n_0_0_5), .ZN(n_0_0_6));
   OAI21_X1 i_0_0_73 (.A(n_0_0_3), .B1(n_0_0_4), .B2(n_0_0_6), .ZN(n_0_128));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_6), .A2(i[3]), .ZN(n_0_0_7));
   OAI211_X1 i_0_0_75 (.A(n_0_0_7), .B(n_0_0_0), .C1(i[3]), .C2(n_0_0_6), 
      .ZN(n_0_0_8));
   NAND2_X1 i_0_0_76 (.A1(start_i[3]), .A2(start), .ZN(n_0_0_9));
   NAND2_X1 i_0_0_77 (.A1(n_0_0_8), .A2(n_0_0_9), .ZN(n_0_129));
   NAND2_X1 i_0_0_78 (.A1(start_i[4]), .A2(start), .ZN(n_0_0_10));
   INV_X1 i_0_0_79 (.A(n_0_0_7), .ZN(n_0_0_11));
   NAND2_X1 i_0_0_80 (.A1(i[4]), .A2(i[3]), .ZN(n_0_0_12));
   OAI22_X1 i_0_0_81 (.A1(n_0_0_11), .A2(i[4]), .B1(n_0_0_5), .B2(n_0_0_12), 
      .ZN(n_0_0_13));
   OAI21_X1 i_0_0_82 (.A(n_0_0_10), .B1(n_0_0_13), .B2(start), .ZN(n_0_130));
   INV_X1 i_0_0_83 (.A(i[3]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_14), .A2(i[4]), .ZN(n_0_0_15));
   INV_X1 i_0_0_85 (.A(i[0]), .ZN(n_0_0_16));
   NOR4_X1 i_0_0_86 (.A1(n_0_0_15), .A2(n_0_0_16), .A3(i[2]), .A4(i[1]), 
      .ZN(n_0_0_17));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_17), .A2(n_0_0_0), .ZN(n_0_131));
   INV_X1 i_0_0_88 (.A(i[1]), .ZN(n_0_0_18));
   INV_X1 i_0_0_89 (.A(n_0_0_12), .ZN(n_0_0_19));
   INV_X1 i_0_0_90 (.A(n_0_0_15), .ZN(n_0_0_20));
   AOI22_X1 i_0_0_91 (.A1(n_0_0_19), .A2(read_data[27]), .B1(n_0_0_20), .B2(
      read_data[19]), .ZN(n_0_0_21));
   OAI22_X1 i_0_0_92 (.A1(n_0_0_14), .A2(read_data[11]), .B1(read_data[3]), 
      .B2(i[3]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_93 (.A(n_0_0_21), .B1(i[4]), .B2(n_0_0_22), .ZN(n_0_0_23));
   INV_X1 i_0_0_94 (.A(n_0_0_23), .ZN(n_0_0_24));
   INV_X1 i_0_0_95 (.A(i[2]), .ZN(n_0_0_25));
   INV_X1 i_0_0_96 (.A(i[4]), .ZN(n_0_0_26));
   AND3_X1 i_0_0_97 (.A1(n_0_0_26), .A2(i[3]), .A3(read_data[7]), .ZN(n_0_0_27));
   AOI221_X1 i_0_0_98 (.A(n_0_0_27), .B1(n_0_0_19), .B2(read_data[23]), .C1(
      read_data[15]), .C2(n_0_0_20), .ZN(n_0_0_28));
   OAI221_X1 i_0_0_99 (.A(n_0_0_18), .B1(n_0_0_24), .B2(n_0_0_25), .C1(n_0_0_28), 
      .C2(i[2]), .ZN(n_0_0_29));
   NOR2_X1 i_0_0_100 (.A1(n_0_0_25), .A2(i[4]), .ZN(n_0_0_30));
   NAND3_X1 i_0_0_101 (.A1(n_0_0_30), .A2(read_data[5]), .A3(n_0_0_14), .ZN(
      n_0_0_31));
   AOI22_X1 i_0_0_102 (.A1(read_data[25]), .A2(n_0_0_19), .B1(n_0_0_20), 
      .B2(read_data[17]), .ZN(n_0_0_32));
   OAI22_X1 i_0_0_103 (.A1(n_0_0_14), .A2(read_data[9]), .B1(read_data[1]), 
      .B2(i[3]), .ZN(n_0_0_33));
   OAI21_X1 i_0_0_104 (.A(n_0_0_32), .B1(i[4]), .B2(n_0_0_33), .ZN(n_0_0_34));
   INV_X1 i_0_0_105 (.A(n_0_0_34), .ZN(n_0_0_35));
   AND3_X1 i_0_0_106 (.A1(n_0_0_26), .A2(read_data[13]), .A3(i[3]), .ZN(n_0_0_36));
   AOI221_X1 i_0_0_107 (.A(n_0_0_36), .B1(read_data[21]), .B2(n_0_0_20), 
      .C1(read_data[29]), .C2(n_0_0_19), .ZN(n_0_0_37));
   OAI221_X1 i_0_0_108 (.A(n_0_0_31), .B1(n_0_0_35), .B2(i[2]), .C1(n_0_0_37), 
      .C2(n_0_0_25), .ZN(n_0_0_38));
   OAI21_X1 i_0_0_109 (.A(n_0_0_29), .B1(n_0_0_38), .B2(n_0_0_18), .ZN(n_0_0_39));
   OAI221_X1 i_0_0_110 (.A(n_0_0_19), .B1(read_data[24]), .B2(i[2]), .C1(
      read_data[28]), .C2(n_0_0_25), .ZN(n_0_0_40));
   OAI221_X1 i_0_0_111 (.A(n_0_0_30), .B1(read_data[4]), .B2(i[3]), .C1(n_0_0_14), 
      .C2(read_data[12]), .ZN(n_0_0_41));
   OAI21_X1 i_0_0_112 (.A(n_0_0_25), .B1(n_0_0_14), .B2(read_data[8]), .ZN(
      n_0_0_42));
   OAI21_X1 i_0_0_113 (.A(n_0_0_26), .B1(read_data[0]), .B2(i[3]), .ZN(n_0_0_43));
   OAI211_X1 i_0_0_114 (.A(n_0_0_40), .B(n_0_0_41), .C1(n_0_0_42), .C2(n_0_0_43), 
      .ZN(n_0_0_44));
   OAI221_X1 i_0_0_115 (.A(n_0_0_20), .B1(read_data[16]), .B2(i[2]), .C1(
      n_0_0_25), .C2(read_data[20]), .ZN(n_0_0_45));
   INV_X1 i_0_0_116 (.A(n_0_0_45), .ZN(n_0_0_46));
   OR3_X1 i_0_0_117 (.A1(n_0_0_44), .A2(i[1]), .A3(n_0_0_46), .ZN(n_0_0_47));
   AOI221_X1 i_0_0_118 (.A(n_0_0_25), .B1(n_0_0_20), .B2(read_data[22]), 
      .C1(n_0_0_19), .C2(read_data[30]), .ZN(n_0_0_48));
   OAI22_X1 i_0_0_119 (.A1(n_0_0_14), .A2(read_data[10]), .B1(read_data[2]), 
      .B2(i[3]), .ZN(n_0_0_49));
   NOR2_X1 i_0_0_120 (.A1(n_0_0_49), .A2(i[4]), .ZN(n_0_0_50));
   AOI221_X1 i_0_0_121 (.A(n_0_0_50), .B1(read_data[26]), .B2(n_0_0_19), 
      .C1(read_data[18]), .C2(n_0_0_20), .ZN(n_0_0_51));
   AOI21_X1 i_0_0_122 (.A(n_0_0_48), .B1(n_0_0_51), .B2(n_0_0_25), .ZN(n_0_0_52));
   OAI221_X1 i_0_0_123 (.A(n_0_0_30), .B1(read_data[6]), .B2(i[3]), .C1(n_0_0_14), 
      .C2(read_data[14]), .ZN(n_0_0_53));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_53), .A2(i[1]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_125 (.A(n_0_0_47), .B1(n_0_0_52), .B2(n_0_0_54), .ZN(n_0_0_55));
   OAI22_X1 i_0_0_126 (.A1(n_0_0_39), .A2(i[0]), .B1(n_0_0_55), .B2(n_0_0_16), 
      .ZN(n_0_0_56));
   OR3_X1 i_0_0_127 (.A1(n_0_0_44), .A2(n_0_0_18), .A3(n_0_0_46), .ZN(n_0_0_57));
   AND3_X1 i_0_0_128 (.A1(n_0_0_26), .A2(read_data[6]), .A3(i[3]), .ZN(n_0_0_58));
   AOI221_X1 i_0_0_129 (.A(n_0_0_58), .B1(n_0_0_19), .B2(read_data[22]), 
      .C1(read_data[14]), .C2(n_0_0_20), .ZN(n_0_0_59));
   AOI22_X1 i_0_0_130 (.A1(n_0_0_51), .A2(i[2]), .B1(n_0_0_59), .B2(n_0_0_25), 
      .ZN(n_0_0_60));
   OAI21_X1 i_0_0_131 (.A(n_0_0_57), .B1(n_0_0_60), .B2(i[1]), .ZN(n_0_0_61));
   AOI22_X1 i_0_0_132 (.A1(n_0_0_39), .A2(i[0]), .B1(n_0_0_61), .B2(n_0_0_16), 
      .ZN(n_0_0_62));
   OR2_X1 i_0_0_133 (.A1(n_0_0_56), .A2(n_0_0_62), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_134 (.A1(n_0_0_56), .A2(n_0_0_62), .ZN(n_0_0_64));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_63), .A2(n_0_0_64), .ZN(n_0_0_65));
   INV_X1 i_0_0_136 (.A(n_0_0_65), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_66), .A2(read_data2[0]), .ZN(n_0_0_67));
   NOR2_X1 i_0_0_138 (.A1(n_0_0_17), .A2(start), .ZN(n_0_0_68));
   INV_X1 i_0_0_139 (.A(shift[4]), .ZN(n_0_0_69));
   INV_X1 i_0_0_140 (.A(shift[2]), .ZN(n_0_0_70));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_69), .A2(n_0_0_70), .ZN(n_0_0_71));
   OR2_X1 i_0_0_142 (.A1(n_0_0_71), .A2(shift[3]), .ZN(n_0_0_72));
   NOR2_X1 i_0_0_143 (.A1(n_0_0_72), .A2(shift[1]), .ZN(n_0_0_73));
   AND2_X1 i_0_0_144 (.A1(n_0_0_68), .A2(n_0_0_73), .ZN(n_0_0_74));
   INV_X1 i_0_0_145 (.A(n_0_0_74), .ZN(n_0_0_75));
   NOR3_X1 i_0_0_146 (.A1(n_0_0_67), .A2(shift[0]), .A3(n_0_0_75), .ZN(n_0_176));
   OAI221_X1 i_0_0_147 (.A(n_0_0_30), .B1(i[3]), .B2(read_data[7]), .C1(n_0_0_14), 
      .C2(read_data[15]), .ZN(n_0_0_76));
   AOI22_X1 i_0_0_148 (.A1(n_0_0_19), .A2(read_data[31]), .B1(n_0_0_20), 
      .B2(read_data[23]), .ZN(n_0_0_77));
   OAI21_X1 i_0_0_149 (.A(n_0_0_76), .B1(n_0_0_25), .B2(n_0_0_77), .ZN(n_0_0_78));
   AOI21_X1 i_0_0_150 (.A(n_0_0_78), .B1(n_0_0_25), .B2(n_0_0_23), .ZN(n_0_0_79));
   INV_X1 i_0_0_151 (.A(n_0_0_38), .ZN(n_0_0_80));
   AOI221_X1 i_0_0_152 (.A(n_0_0_16), .B1(n_0_0_79), .B2(i[1]), .C1(n_0_0_80), 
      .C2(n_0_0_18), .ZN(n_0_0_81));
   INV_X1 i_0_0_153 (.A(n_0_0_55), .ZN(n_0_0_82));
   AOI21_X1 i_0_0_154 (.A(n_0_0_81), .B1(n_0_0_16), .B2(n_0_0_82), .ZN(n_0_0_83));
   INV_X1 i_0_0_155 (.A(n_0_0_83), .ZN(n_0_0_84));
   AND3_X1 i_0_0_156 (.A1(n_0_0_84), .A2(n_0_0_64), .A3(n_0_0_63), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_157 (.A1(n_0_0_65), .A2(n_0_0_84), .ZN(n_0_0_86));
   AOI22_X1 i_0_0_158 (.A1(n_0_0_85), .A2(n_0_9), .B1(n_0_0_86), .B2(
      read_data2[1]), .ZN(n_0_0_87));
   NOR2_X1 i_0_0_159 (.A1(n_0_0_63), .A2(n_0_0_83), .ZN(n_0_0_88));
   NOR2_X1 i_0_0_160 (.A1(n_0_0_84), .A2(n_0_0_64), .ZN(n_0_0_89));
   OAI21_X1 i_0_0_161 (.A(read_data2[0]), .B1(n_0_0_88), .B2(n_0_0_89), .ZN(
      n_0_0_90));
   NAND2_X1 i_0_0_162 (.A1(n_0_0_87), .A2(n_0_0_90), .ZN(n_0_0_91));
   INV_X1 i_0_0_163 (.A(n_0_0_91), .ZN(n_0_0_92));
   INV_X1 i_0_0_164 (.A(shift[0]), .ZN(n_0_0_93));
   AOI221_X1 i_0_0_165 (.A(n_0_0_75), .B1(shift[0]), .B2(n_0_0_67), .C1(n_0_0_92), 
      .C2(n_0_0_93), .ZN(n_0_177));
   INV_X1 i_0_0_166 (.A(n_0_0_68), .ZN(n_0_0_94));
   NOR2_X1 i_0_0_167 (.A1(n_0_0_94), .A2(shift[0]), .ZN(n_0_0_95));
   AOI21_X1 i_0_0_168 (.A(n_0_0_95), .B1(n_0_0_91), .B2(n_0_0_74), .ZN(n_0_0_96));
   AOI22_X1 i_0_0_169 (.A1(n_0_0_85), .A2(n_0_10), .B1(n_0_0_86), .B2(
      read_data2[2]), .ZN(n_0_0_97));
   AOI22_X1 i_0_0_170 (.A1(n_0_0_88), .A2(n_0_40), .B1(n_0_0_89), .B2(
      read_data2[1]), .ZN(n_0_0_98));
   NAND2_X1 i_0_0_171 (.A1(n_0_0_97), .A2(n_0_0_98), .ZN(n_0_0_99));
   INV_X1 i_0_0_172 (.A(n_0_0_67), .ZN(n_0_0_100));
   INV_X1 i_0_0_173 (.A(shift[1]), .ZN(n_0_0_101));
   NOR2_X1 i_0_0_174 (.A1(n_0_0_72), .A2(n_0_0_101), .ZN(n_0_0_102));
   AOI22_X1 i_0_0_175 (.A1(n_0_0_99), .A2(n_0_0_73), .B1(n_0_0_100), .B2(
      n_0_0_102), .ZN(n_0_0_103));
   AOI21_X1 i_0_0_176 (.A(n_0_0_96), .B1(n_0_0_103), .B2(n_0_0_93), .ZN(n_0_178));
   AOI22_X1 i_0_0_177 (.A1(n_0_0_85), .A2(n_0_11), .B1(n_0_0_86), .B2(
      read_data2[3]), .ZN(n_0_0_104));
   AOI22_X1 i_0_0_178 (.A1(n_0_0_88), .A2(n_0_41), .B1(n_0_0_89), .B2(
      read_data2[2]), .ZN(n_0_0_105));
   NAND2_X1 i_0_0_179 (.A1(n_0_0_104), .A2(n_0_0_105), .ZN(n_0_0_106));
   AOI22_X1 i_0_0_180 (.A1(n_0_0_91), .A2(n_0_0_102), .B1(n_0_0_106), .B2(
      n_0_0_73), .ZN(n_0_0_107));
   INV_X1 i_0_0_181 (.A(n_0_0_95), .ZN(n_0_0_108));
   NAND2_X1 i_0_0_182 (.A1(n_0_0_68), .A2(shift[0]), .ZN(n_0_0_109));
   OAI22_X1 i_0_0_183 (.A1(n_0_0_107), .A2(n_0_0_108), .B1(n_0_0_103), .B2(
      n_0_0_109), .ZN(n_0_179));
   AOI22_X1 i_0_0_184 (.A1(n_0_0_85), .A2(n_0_12), .B1(n_0_0_86), .B2(
      read_data2[4]), .ZN(n_0_0_110));
   AOI22_X1 i_0_0_185 (.A1(n_0_0_88), .A2(n_0_42), .B1(n_0_0_89), .B2(
      read_data2[3]), .ZN(n_0_0_111));
   NAND2_X1 i_0_0_186 (.A1(n_0_0_110), .A2(n_0_0_111), .ZN(n_0_0_112));
   INV_X1 i_0_0_187 (.A(n_0_0_112), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_69), .A2(shift[2]), .ZN(n_0_0_114));
   OR2_X1 i_0_0_189 (.A1(n_0_0_114), .A2(shift[3]), .ZN(n_0_0_115));
   OAI22_X1 i_0_0_190 (.A1(n_0_0_113), .A2(n_0_0_72), .B1(n_0_0_67), .B2(
      n_0_0_115), .ZN(n_0_0_116));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_116), .A2(n_0_0_101), .B1(n_0_0_99), .B2(
      n_0_0_102), .ZN(n_0_0_117));
   OAI22_X1 i_0_0_192 (.A1(n_0_0_117), .A2(n_0_0_108), .B1(n_0_0_109), .B2(
      n_0_0_107), .ZN(n_0_180));
   AOI22_X1 i_0_0_193 (.A1(n_0_0_85), .A2(n_0_13), .B1(n_0_0_86), .B2(
      read_data2[5]), .ZN(n_0_0_118));
   AOI22_X1 i_0_0_194 (.A1(n_0_0_88), .A2(n_0_43), .B1(n_0_0_89), .B2(
      read_data2[4]), .ZN(n_0_0_119));
   NAND2_X1 i_0_0_195 (.A1(n_0_0_118), .A2(n_0_0_119), .ZN(n_0_0_120));
   INV_X1 i_0_0_196 (.A(n_0_0_120), .ZN(n_0_0_121));
   OAI22_X1 i_0_0_197 (.A1(n_0_0_121), .A2(n_0_0_72), .B1(n_0_0_92), .B2(
      n_0_0_115), .ZN(n_0_0_122));
   AOI22_X1 i_0_0_198 (.A1(n_0_0_122), .A2(n_0_0_101), .B1(n_0_0_106), .B2(
      n_0_0_102), .ZN(n_0_0_123));
   OAI22_X1 i_0_0_199 (.A1(n_0_0_123), .A2(n_0_0_108), .B1(n_0_0_117), .B2(
      n_0_0_109), .ZN(n_0_181));
   INV_X1 i_0_0_200 (.A(n_0_0_99), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_201 (.A1(n_0_0_85), .A2(n_0_14), .B1(n_0_0_86), .B2(
      read_data2[6]), .ZN(n_0_0_125));
   AOI22_X1 i_0_0_202 (.A1(n_0_0_88), .A2(n_0_44), .B1(n_0_0_89), .B2(
      read_data2[5]), .ZN(n_0_0_126));
   NAND2_X1 i_0_0_203 (.A1(n_0_0_125), .A2(n_0_0_126), .ZN(n_0_0_127));
   INV_X1 i_0_0_204 (.A(n_0_0_127), .ZN(n_0_0_128));
   OAI22_X1 i_0_0_205 (.A1(n_0_0_124), .A2(n_0_0_115), .B1(n_0_0_128), .B2(
      n_0_0_72), .ZN(n_0_0_129));
   AOI22_X1 i_0_0_206 (.A1(n_0_0_129), .A2(n_0_0_101), .B1(n_0_0_116), .B2(
      shift[1]), .ZN(n_0_0_130));
   OAI22_X1 i_0_0_207 (.A1(n_0_0_130), .A2(n_0_0_108), .B1(n_0_0_123), .B2(
      n_0_0_109), .ZN(n_0_182));
   AOI22_X1 i_0_0_208 (.A1(n_0_0_85), .A2(n_0_15), .B1(n_0_0_86), .B2(
      read_data2[7]), .ZN(n_0_0_131));
   AOI22_X1 i_0_0_209 (.A1(n_0_0_88), .A2(n_0_45), .B1(n_0_0_89), .B2(
      read_data2[6]), .ZN(n_0_0_132));
   NAND2_X1 i_0_0_210 (.A1(n_0_0_131), .A2(n_0_0_132), .ZN(n_0_0_133));
   INV_X1 i_0_0_211 (.A(n_0_0_133), .ZN(n_0_0_134));
   INV_X1 i_0_0_212 (.A(n_0_0_106), .ZN(n_0_0_135));
   OAI22_X1 i_0_0_213 (.A1(n_0_0_134), .A2(n_0_0_72), .B1(n_0_0_135), .B2(
      n_0_0_115), .ZN(n_0_0_136));
   AOI22_X1 i_0_0_214 (.A1(n_0_0_122), .A2(shift[1]), .B1(n_0_0_136), .B2(
      n_0_0_101), .ZN(n_0_0_137));
   OAI22_X1 i_0_0_215 (.A1(n_0_0_137), .A2(n_0_0_108), .B1(n_0_0_130), .B2(
      n_0_0_109), .ZN(n_0_183));
   AOI22_X1 i_0_0_216 (.A1(n_0_0_85), .A2(n_0_16), .B1(n_0_0_86), .B2(
      read_data2[8]), .ZN(n_0_0_138));
   AOI22_X1 i_0_0_217 (.A1(n_0_0_88), .A2(n_0_46), .B1(n_0_0_89), .B2(
      read_data2[7]), .ZN(n_0_0_139));
   NAND2_X1 i_0_0_218 (.A1(n_0_0_138), .A2(n_0_0_139), .ZN(n_0_0_140));
   NOR2_X1 i_0_0_219 (.A1(shift[4]), .A2(shift[3]), .ZN(n_0_0_141));
   INV_X1 i_0_0_220 (.A(shift[3]), .ZN(n_0_0_142));
   NOR2_X1 i_0_0_221 (.A1(n_0_0_142), .A2(shift[4]), .ZN(n_0_0_143));
   AOI22_X1 i_0_0_222 (.A1(n_0_0_140), .A2(n_0_0_141), .B1(n_0_0_100), .B2(
      n_0_0_143), .ZN(n_0_0_144));
   OAI22_X1 i_0_0_223 (.A1(n_0_0_144), .A2(shift[2]), .B1(n_0_0_113), .B2(
      n_0_0_115), .ZN(n_0_0_145));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_145), .A2(n_0_0_101), .B1(n_0_0_129), .B2(
      shift[1]), .ZN(n_0_0_146));
   OAI22_X1 i_0_0_225 (.A1(n_0_0_146), .A2(n_0_0_108), .B1(n_0_0_137), .B2(
      n_0_0_109), .ZN(n_0_184));
   AOI22_X1 i_0_0_226 (.A1(n_0_0_85), .A2(n_0_17), .B1(n_0_0_86), .B2(
      read_data2[9]), .ZN(n_0_0_147));
   AOI22_X1 i_0_0_227 (.A1(n_0_0_88), .A2(n_0_47), .B1(n_0_0_89), .B2(
      read_data2[8]), .ZN(n_0_0_148));
   NAND2_X1 i_0_0_228 (.A1(n_0_0_147), .A2(n_0_0_148), .ZN(n_0_0_149));
   AOI22_X1 i_0_0_229 (.A1(n_0_0_91), .A2(n_0_0_143), .B1(n_0_0_149), .B2(
      n_0_0_141), .ZN(n_0_0_150));
   OAI22_X1 i_0_0_230 (.A1(n_0_0_150), .A2(shift[2]), .B1(n_0_0_121), .B2(
      n_0_0_115), .ZN(n_0_0_151));
   AOI22_X1 i_0_0_231 (.A1(n_0_0_151), .A2(n_0_0_101), .B1(n_0_0_136), .B2(
      shift[1]), .ZN(n_0_0_152));
   OAI22_X1 i_0_0_232 (.A1(n_0_0_152), .A2(n_0_0_108), .B1(n_0_0_146), .B2(
      n_0_0_109), .ZN(n_0_185));
   AOI22_X1 i_0_0_233 (.A1(n_0_0_85), .A2(n_0_18), .B1(n_0_0_86), .B2(
      read_data2[10]), .ZN(n_0_0_153));
   AOI22_X1 i_0_0_234 (.A1(n_0_0_88), .A2(n_0_48), .B1(n_0_0_89), .B2(
      read_data2[9]), .ZN(n_0_0_154));
   NAND2_X1 i_0_0_235 (.A1(n_0_0_153), .A2(n_0_0_154), .ZN(n_0_0_155));
   AOI22_X1 i_0_0_236 (.A1(n_0_0_99), .A2(shift[3]), .B1(n_0_0_155), .B2(
      n_0_0_142), .ZN(n_0_0_156));
   OAI22_X1 i_0_0_237 (.A1(n_0_0_156), .A2(n_0_0_71), .B1(n_0_0_128), .B2(
      n_0_0_115), .ZN(n_0_0_157));
   AOI22_X1 i_0_0_238 (.A1(n_0_0_157), .A2(n_0_0_101), .B1(n_0_0_145), .B2(
      shift[1]), .ZN(n_0_0_158));
   OAI22_X1 i_0_0_239 (.A1(n_0_0_152), .A2(n_0_0_109), .B1(n_0_0_158), .B2(
      n_0_0_108), .ZN(n_0_186));
   AOI22_X1 i_0_0_240 (.A1(n_0_0_85), .A2(n_0_19), .B1(n_0_0_86), .B2(
      read_data2[11]), .ZN(n_0_0_159));
   AOI22_X1 i_0_0_241 (.A1(n_0_0_88), .A2(n_0_49), .B1(n_0_0_89), .B2(
      read_data2[10]), .ZN(n_0_0_160));
   NAND2_X1 i_0_0_242 (.A1(n_0_0_159), .A2(n_0_0_160), .ZN(n_0_0_161));
   AOI22_X1 i_0_0_243 (.A1(n_0_0_161), .A2(n_0_0_142), .B1(n_0_0_106), .B2(
      shift[3]), .ZN(n_0_0_162));
   OAI22_X1 i_0_0_244 (.A1(n_0_0_162), .A2(n_0_0_71), .B1(n_0_0_134), .B2(
      n_0_0_115), .ZN(n_0_0_163));
   AOI22_X1 i_0_0_245 (.A1(n_0_0_163), .A2(n_0_0_101), .B1(n_0_0_151), .B2(
      shift[1]), .ZN(n_0_0_164));
   OAI22_X1 i_0_0_246 (.A1(n_0_0_164), .A2(n_0_0_108), .B1(n_0_0_158), .B2(
      n_0_0_109), .ZN(n_0_187));
   AOI22_X1 i_0_0_247 (.A1(n_0_0_85), .A2(n_0_20), .B1(n_0_0_86), .B2(
      read_data2[12]), .ZN(n_0_0_165));
   AOI22_X1 i_0_0_248 (.A1(n_0_0_88), .A2(n_0_50), .B1(n_0_0_89), .B2(
      read_data2[11]), .ZN(n_0_0_166));
   NAND2_X1 i_0_0_249 (.A1(n_0_0_165), .A2(n_0_0_166), .ZN(n_0_0_167));
   AOI22_X1 i_0_0_250 (.A1(n_0_0_167), .A2(n_0_0_142), .B1(n_0_0_112), .B2(
      shift[3]), .ZN(n_0_0_168));
   OAI22_X1 i_0_0_251 (.A1(n_0_0_168), .A2(n_0_0_71), .B1(n_0_0_144), .B2(
      n_0_0_70), .ZN(n_0_0_169));
   AOI22_X1 i_0_0_252 (.A1(n_0_0_101), .A2(n_0_0_169), .B1(n_0_0_157), .B2(
      shift[1]), .ZN(n_0_0_170));
   OAI22_X1 i_0_0_253 (.A1(n_0_0_164), .A2(n_0_0_109), .B1(n_0_0_170), .B2(
      n_0_0_108), .ZN(n_0_188));
   AOI22_X1 i_0_0_254 (.A1(n_0_0_85), .A2(n_0_21), .B1(n_0_0_86), .B2(
      read_data2[13]), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_255 (.A1(n_0_0_88), .A2(n_0_51), .B1(n_0_0_89), .B2(
      read_data2[12]), .ZN(n_0_0_172));
   NAND2_X1 i_0_0_256 (.A1(n_0_0_171), .A2(n_0_0_172), .ZN(n_0_0_173));
   AOI22_X1 i_0_0_257 (.A1(n_0_0_120), .A2(shift[3]), .B1(n_0_0_173), .B2(
      n_0_0_142), .ZN(n_0_0_174));
   OAI22_X1 i_0_0_258 (.A1(n_0_0_150), .A2(n_0_0_70), .B1(n_0_0_174), .B2(
      n_0_0_71), .ZN(n_0_0_175));
   AOI22_X1 i_0_0_259 (.A1(n_0_0_175), .A2(n_0_0_101), .B1(n_0_0_163), .B2(
      shift[1]), .ZN(n_0_0_176));
   OAI22_X1 i_0_0_260 (.A1(n_0_0_176), .A2(n_0_0_108), .B1(n_0_0_170), .B2(
      n_0_0_109), .ZN(n_0_189));
   AOI22_X1 i_0_0_261 (.A1(n_0_0_85), .A2(n_0_22), .B1(n_0_0_86), .B2(
      read_data2[14]), .ZN(n_0_0_177));
   AOI22_X1 i_0_0_262 (.A1(n_0_0_88), .A2(n_0_52), .B1(n_0_0_89), .B2(
      read_data2[13]), .ZN(n_0_0_178));
   NAND2_X1 i_0_0_263 (.A1(n_0_0_177), .A2(n_0_0_178), .ZN(n_0_0_179));
   AOI22_X1 i_0_0_264 (.A1(n_0_0_179), .A2(n_0_0_141), .B1(n_0_0_127), .B2(
      n_0_0_143), .ZN(n_0_0_180));
   OAI22_X1 i_0_0_265 (.A1(n_0_0_156), .A2(n_0_0_114), .B1(n_0_0_180), .B2(
      shift[2]), .ZN(n_0_0_181));
   AOI22_X1 i_0_0_266 (.A1(n_0_0_181), .A2(n_0_0_101), .B1(n_0_0_169), .B2(
      shift[1]), .ZN(n_0_0_182));
   OAI22_X1 i_0_0_267 (.A1(n_0_0_176), .A2(n_0_0_109), .B1(n_0_0_182), .B2(
      n_0_0_108), .ZN(n_0_190));
   AOI22_X1 i_0_0_268 (.A1(n_0_0_85), .A2(n_0_23), .B1(n_0_0_86), .B2(
      read_data2[15]), .ZN(n_0_0_183));
   AOI22_X1 i_0_0_269 (.A1(n_0_0_88), .A2(n_0_53), .B1(n_0_0_89), .B2(
      read_data2[14]), .ZN(n_0_0_184));
   NAND2_X1 i_0_0_270 (.A1(n_0_0_183), .A2(n_0_0_184), .ZN(n_0_0_185));
   AOI22_X1 i_0_0_271 (.A1(n_0_0_133), .A2(shift[3]), .B1(n_0_0_185), .B2(
      n_0_0_142), .ZN(n_0_0_186));
   OAI22_X1 i_0_0_272 (.A1(n_0_0_162), .A2(n_0_0_114), .B1(n_0_0_186), .B2(
      n_0_0_71), .ZN(n_0_0_187));
   AOI22_X1 i_0_0_273 (.A1(n_0_0_175), .A2(shift[1]), .B1(n_0_0_187), .B2(
      n_0_0_101), .ZN(n_0_0_188));
   OAI22_X1 i_0_0_274 (.A1(n_0_0_188), .A2(n_0_0_108), .B1(n_0_0_182), .B2(
      n_0_0_109), .ZN(n_0_191));
   AOI22_X1 i_0_0_275 (.A1(n_0_0_85), .A2(n_0_24), .B1(n_0_0_86), .B2(
      read_data2[16]), .ZN(n_0_0_189));
   AOI22_X1 i_0_0_276 (.A1(n_0_0_88), .A2(n_0_54), .B1(n_0_0_89), .B2(
      read_data2[15]), .ZN(n_0_0_190));
   NAND2_X1 i_0_0_277 (.A1(n_0_0_189), .A2(n_0_0_190), .ZN(n_0_0_191));
   INV_X1 i_0_0_278 (.A(n_0_0_191), .ZN(n_0_0_192));
   AOI22_X1 i_0_0_279 (.A1(n_0_0_192), .A2(n_0_0_69), .B1(n_0_0_67), .B2(
      shift[4]), .ZN(n_0_0_193));
   AOI22_X1 i_0_0_280 (.A1(n_0_0_193), .A2(n_0_0_142), .B1(n_0_0_140), .B2(
      n_0_0_143), .ZN(n_0_0_194));
   OAI22_X1 i_0_0_281 (.A1(n_0_0_194), .A2(shift[2]), .B1(n_0_0_168), .B2(
      n_0_0_114), .ZN(n_0_0_195));
   AOI22_X1 i_0_0_282 (.A1(n_0_0_195), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_181), .ZN(n_0_0_196));
   OAI22_X1 i_0_0_283 (.A1(n_0_0_196), .A2(n_0_0_108), .B1(n_0_0_188), .B2(
      n_0_0_109), .ZN(n_0_192));
   AOI22_X1 i_0_0_284 (.A1(n_0_0_85), .A2(n_0_25), .B1(n_0_0_86), .B2(
      read_data2[17]), .ZN(n_0_0_197));
   AOI22_X1 i_0_0_285 (.A1(n_0_0_88), .A2(n_0_55), .B1(n_0_0_89), .B2(
      read_data2[16]), .ZN(n_0_0_198));
   NAND2_X1 i_0_0_286 (.A1(n_0_0_197), .A2(n_0_0_198), .ZN(n_0_0_199));
   INV_X1 i_0_0_287 (.A(n_0_0_199), .ZN(n_0_0_200));
   OAI22_X1 i_0_0_288 (.A1(n_0_0_200), .A2(shift[4]), .B1(n_0_0_92), .B2(
      n_0_0_69), .ZN(n_0_0_201));
   AOI22_X1 i_0_0_289 (.A1(n_0_0_201), .A2(n_0_0_142), .B1(n_0_0_149), .B2(
      n_0_0_143), .ZN(n_0_0_202));
   OAI22_X1 i_0_0_290 (.A1(n_0_0_202), .A2(shift[2]), .B1(n_0_0_174), .B2(
      n_0_0_114), .ZN(n_0_0_203));
   INV_X1 i_0_0_291 (.A(n_0_0_203), .ZN(n_0_0_204));
   INV_X1 i_0_0_292 (.A(n_0_0_187), .ZN(n_0_0_205));
   AOI22_X1 i_0_0_293 (.A1(n_0_0_204), .A2(n_0_0_101), .B1(n_0_0_205), .B2(
      shift[1]), .ZN(n_0_0_206));
   NAND2_X1 i_0_0_294 (.A1(n_0_0_206), .A2(n_0_0_68), .ZN(n_0_0_207));
   AOI22_X1 i_0_0_295 (.A1(n_0_0_207), .A2(n_0_0_109), .B1(shift[0]), .B2(
      n_0_0_196), .ZN(n_0_193));
   AOI22_X1 i_0_0_296 (.A1(n_0_0_85), .A2(n_0_26), .B1(n_0_0_86), .B2(
      read_data2[18]), .ZN(n_0_0_208));
   AOI22_X1 i_0_0_297 (.A1(n_0_0_88), .A2(n_0_56), .B1(n_0_0_89), .B2(
      read_data2[17]), .ZN(n_0_0_209));
   NAND2_X1 i_0_0_298 (.A1(n_0_0_208), .A2(n_0_0_209), .ZN(n_0_0_210));
   INV_X1 i_0_0_299 (.A(n_0_0_210), .ZN(n_0_0_211));
   OAI22_X1 i_0_0_300 (.A1(n_0_0_211), .A2(shift[4]), .B1(n_0_0_124), .B2(
      n_0_0_69), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_301 (.A1(n_0_0_212), .A2(n_0_0_142), .B1(n_0_0_155), .B2(
      n_0_0_143), .ZN(n_0_0_213));
   OAI22_X1 i_0_0_302 (.A1(n_0_0_213), .A2(shift[2]), .B1(n_0_0_70), .B2(
      n_0_0_180), .ZN(n_0_0_214));
   AOI22_X1 i_0_0_303 (.A1(n_0_0_214), .A2(n_0_0_101), .B1(n_0_0_195), .B2(
      shift[1]), .ZN(n_0_0_215));
   AOI22_X1 i_0_0_304 (.A1(n_0_0_207), .A2(n_0_0_108), .B1(n_0_0_215), .B2(
      n_0_0_93), .ZN(n_0_194));
   AOI22_X1 i_0_0_305 (.A1(n_0_0_85), .A2(n_0_27), .B1(n_0_0_86), .B2(
      read_data2[19]), .ZN(n_0_0_216));
   AOI22_X1 i_0_0_306 (.A1(n_0_0_88), .A2(n_0_57), .B1(n_0_0_89), .B2(
      read_data2[18]), .ZN(n_0_0_217));
   NAND2_X1 i_0_0_307 (.A1(n_0_0_216), .A2(n_0_0_217), .ZN(n_0_0_218));
   INV_X1 i_0_0_308 (.A(n_0_0_218), .ZN(n_0_0_219));
   OAI22_X1 i_0_0_309 (.A1(n_0_0_135), .A2(n_0_0_69), .B1(n_0_0_219), .B2(
      shift[4]), .ZN(n_0_0_220));
   AOI22_X1 i_0_0_310 (.A1(n_0_0_220), .A2(n_0_0_142), .B1(n_0_0_161), .B2(
      n_0_0_143), .ZN(n_0_0_221));
   OAI22_X1 i_0_0_311 (.A1(n_0_0_221), .A2(shift[2]), .B1(n_0_0_186), .B2(
      n_0_0_114), .ZN(n_0_0_222));
   AOI22_X1 i_0_0_312 (.A1(n_0_0_222), .A2(n_0_0_101), .B1(n_0_0_203), .B2(
      shift[1]), .ZN(n_0_0_223));
   OAI22_X1 i_0_0_313 (.A1(n_0_0_223), .A2(n_0_0_108), .B1(n_0_0_215), .B2(
      n_0_0_109), .ZN(n_0_195));
   AOI22_X1 i_0_0_314 (.A1(n_0_0_85), .A2(n_0_28), .B1(n_0_0_86), .B2(
      read_data2[20]), .ZN(n_0_0_224));
   AOI22_X1 i_0_0_315 (.A1(n_0_0_88), .A2(n_0_58), .B1(n_0_0_89), .B2(
      read_data2[19]), .ZN(n_0_0_225));
   NAND2_X1 i_0_0_316 (.A1(n_0_0_224), .A2(n_0_0_225), .ZN(n_0_0_226));
   INV_X1 i_0_0_317 (.A(n_0_0_226), .ZN(n_0_0_227));
   OAI22_X1 i_0_0_318 (.A1(n_0_0_113), .A2(n_0_0_69), .B1(n_0_0_227), .B2(
      shift[4]), .ZN(n_0_0_228));
   AOI22_X1 i_0_0_319 (.A1(n_0_0_228), .A2(n_0_0_142), .B1(n_0_0_167), .B2(
      n_0_0_143), .ZN(n_0_0_229));
   OAI22_X1 i_0_0_320 (.A1(n_0_0_229), .A2(shift[2]), .B1(n_0_0_194), .B2(
      n_0_0_70), .ZN(n_0_0_230));
   AOI22_X1 i_0_0_321 (.A1(n_0_0_101), .A2(n_0_0_230), .B1(n_0_0_214), .B2(
      shift[1]), .ZN(n_0_0_231));
   OAI22_X1 i_0_0_322 (.A1(n_0_0_223), .A2(n_0_0_109), .B1(n_0_0_231), .B2(
      n_0_0_108), .ZN(n_0_196));
   AOI22_X1 i_0_0_323 (.A1(n_0_0_85), .A2(n_0_29), .B1(n_0_0_86), .B2(
      read_data2[21]), .ZN(n_0_0_232));
   AOI22_X1 i_0_0_324 (.A1(n_0_0_88), .A2(n_0_59), .B1(n_0_0_89), .B2(
      read_data2[20]), .ZN(n_0_0_233));
   AND2_X1 i_0_0_325 (.A1(n_0_0_232), .A2(n_0_0_233), .ZN(n_0_0_234));
   OAI22_X1 i_0_0_326 (.A1(n_0_0_234), .A2(shift[4]), .B1(n_0_0_121), .B2(
      n_0_0_69), .ZN(n_0_0_235));
   AOI22_X1 i_0_0_327 (.A1(n_0_0_235), .A2(n_0_0_142), .B1(n_0_0_173), .B2(
      n_0_0_143), .ZN(n_0_0_236));
   OAI22_X1 i_0_0_328 (.A1(n_0_0_236), .A2(shift[2]), .B1(n_0_0_202), .B2(
      n_0_0_70), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_329 (.A1(n_0_0_237), .A2(n_0_0_101), .B1(n_0_0_222), .B2(
      shift[1]), .ZN(n_0_0_238));
   OAI22_X1 i_0_0_330 (.A1(n_0_0_238), .A2(n_0_0_108), .B1(n_0_0_231), .B2(
      n_0_0_109), .ZN(n_0_197));
   AOI22_X1 i_0_0_331 (.A1(n_0_0_85), .A2(n_0_30), .B1(n_0_0_86), .B2(
      read_data2[22]), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_332 (.A1(n_0_0_88), .A2(n_0_60), .B1(n_0_0_89), .B2(
      read_data2[21]), .ZN(n_0_0_240));
   AND2_X1 i_0_0_333 (.A1(n_0_0_239), .A2(n_0_0_240), .ZN(n_0_0_241));
   OAI22_X1 i_0_0_334 (.A1(n_0_0_241), .A2(shift[4]), .B1(n_0_0_128), .B2(
      n_0_0_69), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_335 (.A1(n_0_0_242), .A2(n_0_0_142), .B1(n_0_0_179), .B2(
      n_0_0_143), .ZN(n_0_0_243));
   OAI22_X1 i_0_0_336 (.A1(n_0_0_243), .A2(shift[2]), .B1(n_0_0_213), .B2(
      n_0_0_70), .ZN(n_0_0_244));
   AOI22_X1 i_0_0_337 (.A1(n_0_0_244), .A2(n_0_0_101), .B1(n_0_0_230), .B2(
      shift[1]), .ZN(n_0_0_245));
   OAI22_X1 i_0_0_338 (.A1(n_0_0_245), .A2(n_0_0_108), .B1(n_0_0_238), .B2(
      n_0_0_109), .ZN(n_0_198));
   AOI22_X1 i_0_0_339 (.A1(n_0_0_85), .A2(n_0_31), .B1(n_0_0_86), .B2(
      read_data2[23]), .ZN(n_0_0_246));
   AOI22_X1 i_0_0_340 (.A1(n_0_0_88), .A2(n_0_61), .B1(n_0_0_89), .B2(
      read_data2[22]), .ZN(n_0_0_247));
   AND2_X1 i_0_0_341 (.A1(n_0_0_246), .A2(n_0_0_247), .ZN(n_0_0_248));
   OAI22_X1 i_0_0_342 (.A1(n_0_0_248), .A2(shift[4]), .B1(n_0_0_134), .B2(
      n_0_0_69), .ZN(n_0_0_249));
   AOI22_X1 i_0_0_343 (.A1(n_0_0_249), .A2(n_0_0_142), .B1(n_0_0_185), .B2(
      n_0_0_143), .ZN(n_0_0_250));
   OAI22_X1 i_0_0_344 (.A1(n_0_0_221), .A2(n_0_0_70), .B1(n_0_0_250), .B2(
      shift[2]), .ZN(n_0_0_251));
   AOI22_X1 i_0_0_345 (.A1(n_0_0_237), .A2(shift[1]), .B1(n_0_0_251), .B2(
      n_0_0_101), .ZN(n_0_0_252));
   OAI22_X1 i_0_0_346 (.A1(n_0_0_252), .A2(n_0_0_108), .B1(n_0_0_245), .B2(
      n_0_0_109), .ZN(n_0_199));
   AOI22_X1 i_0_0_347 (.A1(n_0_0_85), .A2(n_0_32), .B1(n_0_0_86), .B2(
      read_data2[24]), .ZN(n_0_0_253));
   AOI22_X1 i_0_0_348 (.A1(n_0_0_88), .A2(n_0_62), .B1(n_0_0_89), .B2(
      read_data2[23]), .ZN(n_0_0_254));
   NAND2_X1 i_0_0_349 (.A1(n_0_0_253), .A2(n_0_0_254), .ZN(n_0_0_255));
   INV_X1 i_0_0_350 (.A(n_0_0_255), .ZN(n_0_0_256));
   INV_X1 i_0_0_351 (.A(n_0_0_140), .ZN(n_0_0_257));
   OAI22_X1 i_0_0_352 (.A1(n_0_0_256), .A2(shift[4]), .B1(n_0_0_257), .B2(
      n_0_0_69), .ZN(n_0_0_258));
   OAI22_X1 i_0_0_353 (.A1(n_0_0_258), .A2(shift[3]), .B1(n_0_0_193), .B2(
      n_0_0_142), .ZN(n_0_0_259));
   OAI22_X1 i_0_0_354 (.A1(n_0_0_259), .A2(shift[2]), .B1(n_0_0_229), .B2(
      n_0_0_70), .ZN(n_0_0_260));
   AOI22_X1 i_0_0_355 (.A1(n_0_0_244), .A2(shift[1]), .B1(n_0_0_260), .B2(
      n_0_0_101), .ZN(n_0_0_261));
   OAI22_X1 i_0_0_356 (.A1(n_0_0_252), .A2(n_0_0_109), .B1(n_0_0_261), .B2(
      n_0_0_108), .ZN(n_0_200));
   INV_X1 i_0_0_357 (.A(n_0_0_149), .ZN(n_0_0_262));
   AOI22_X1 i_0_0_358 (.A1(n_0_0_85), .A2(n_0_33), .B1(n_0_0_86), .B2(
      read_data2[25]), .ZN(n_0_0_263));
   AOI22_X1 i_0_0_359 (.A1(n_0_0_88), .A2(n_0_63), .B1(n_0_0_89), .B2(
      read_data2[24]), .ZN(n_0_0_264));
   NAND2_X1 i_0_0_360 (.A1(n_0_0_263), .A2(n_0_0_264), .ZN(n_0_0_265));
   INV_X1 i_0_0_361 (.A(n_0_0_265), .ZN(n_0_0_266));
   OAI22_X1 i_0_0_362 (.A1(n_0_0_262), .A2(n_0_0_69), .B1(n_0_0_266), .B2(
      shift[4]), .ZN(n_0_0_267));
   AOI22_X1 i_0_0_363 (.A1(n_0_0_201), .A2(shift[3]), .B1(n_0_0_267), .B2(
      n_0_0_142), .ZN(n_0_0_268));
   OAI22_X1 i_0_0_364 (.A1(n_0_0_268), .A2(shift[2]), .B1(n_0_0_236), .B2(
      n_0_0_70), .ZN(n_0_0_269));
   AOI22_X1 i_0_0_365 (.A1(n_0_0_269), .A2(n_0_0_101), .B1(n_0_0_251), .B2(
      shift[1]), .ZN(n_0_0_270));
   OAI22_X1 i_0_0_366 (.A1(n_0_0_270), .A2(n_0_0_108), .B1(n_0_0_261), .B2(
      n_0_0_109), .ZN(n_0_201));
   INV_X1 i_0_0_367 (.A(n_0_0_155), .ZN(n_0_0_271));
   AOI22_X1 i_0_0_368 (.A1(n_0_0_85), .A2(n_0_34), .B1(n_0_0_86), .B2(
      read_data2[26]), .ZN(n_0_0_272));
   AOI22_X1 i_0_0_369 (.A1(n_0_0_88), .A2(n_0_64), .B1(n_0_0_89), .B2(
      read_data2[25]), .ZN(n_0_0_273));
   NAND2_X1 i_0_0_370 (.A1(n_0_0_272), .A2(n_0_0_273), .ZN(n_0_0_274));
   INV_X1 i_0_0_371 (.A(n_0_0_274), .ZN(n_0_0_275));
   OAI22_X1 i_0_0_372 (.A1(n_0_0_271), .A2(n_0_0_69), .B1(n_0_0_275), .B2(
      shift[4]), .ZN(n_0_0_276));
   AOI22_X1 i_0_0_373 (.A1(n_0_0_276), .A2(n_0_0_142), .B1(n_0_0_212), .B2(
      shift[3]), .ZN(n_0_0_277));
   OAI22_X1 i_0_0_374 (.A1(n_0_0_277), .A2(shift[2]), .B1(n_0_0_243), .B2(
      n_0_0_70), .ZN(n_0_0_278));
   AOI22_X1 i_0_0_375 (.A1(n_0_0_278), .A2(n_0_0_101), .B1(n_0_0_260), .B2(
      shift[1]), .ZN(n_0_0_279));
   OAI22_X1 i_0_0_376 (.A1(n_0_0_279), .A2(n_0_0_108), .B1(n_0_0_270), .B2(
      n_0_0_109), .ZN(n_0_132));
   AOI22_X1 i_0_0_377 (.A1(n_0_0_85), .A2(n_0_35), .B1(n_0_0_86), .B2(
      read_data2[27]), .ZN(n_0_0_280));
   AOI22_X1 i_0_0_378 (.A1(n_0_0_88), .A2(n_0_65), .B1(n_0_0_89), .B2(
      read_data2[26]), .ZN(n_0_0_281));
   NAND2_X1 i_0_0_379 (.A1(n_0_0_280), .A2(n_0_0_281), .ZN(n_0_0_282));
   INV_X1 i_0_0_380 (.A(n_0_0_282), .ZN(n_0_0_283));
   INV_X1 i_0_0_381 (.A(n_0_0_161), .ZN(n_0_0_284));
   OAI22_X1 i_0_0_382 (.A1(n_0_0_283), .A2(shift[4]), .B1(n_0_0_284), .B2(
      n_0_0_69), .ZN(n_0_0_285));
   AOI22_X1 i_0_0_383 (.A1(n_0_0_285), .A2(n_0_0_142), .B1(n_0_0_220), .B2(
      shift[3]), .ZN(n_0_0_286));
   OAI22_X1 i_0_0_384 (.A1(n_0_0_286), .A2(shift[2]), .B1(n_0_0_250), .B2(
      n_0_0_70), .ZN(n_0_0_287));
   AOI22_X1 i_0_0_385 (.A1(n_0_0_287), .A2(n_0_0_101), .B1(n_0_0_269), .B2(
      shift[1]), .ZN(n_0_0_288));
   OAI22_X1 i_0_0_386 (.A1(n_0_0_288), .A2(n_0_0_108), .B1(n_0_0_279), .B2(
      n_0_0_109), .ZN(n_0_133));
   INV_X1 i_0_0_387 (.A(n_0_0_167), .ZN(n_0_0_289));
   AOI22_X1 i_0_0_388 (.A1(n_0_0_85), .A2(n_0_36), .B1(n_0_0_86), .B2(
      read_data2[28]), .ZN(n_0_0_290));
   AOI22_X1 i_0_0_389 (.A1(n_0_0_88), .A2(n_0_66), .B1(n_0_0_89), .B2(
      read_data2[27]), .ZN(n_0_0_291));
   AND2_X1 i_0_0_390 (.A1(n_0_0_290), .A2(n_0_0_291), .ZN(n_0_0_292));
   OAI22_X1 i_0_0_391 (.A1(n_0_0_289), .A2(n_0_0_69), .B1(n_0_0_292), .B2(
      shift[4]), .ZN(n_0_0_293));
   AOI22_X1 i_0_0_392 (.A1(n_0_0_293), .A2(n_0_0_142), .B1(n_0_0_228), .B2(
      shift[3]), .ZN(n_0_0_294));
   OAI22_X1 i_0_0_393 (.A1(n_0_0_294), .A2(shift[2]), .B1(n_0_0_259), .B2(
      n_0_0_70), .ZN(n_0_0_295));
   AOI22_X1 i_0_0_394 (.A1(n_0_0_101), .A2(n_0_0_295), .B1(n_0_0_278), .B2(
      shift[1]), .ZN(n_0_0_296));
   OAI22_X1 i_0_0_395 (.A1(n_0_0_288), .A2(n_0_0_109), .B1(n_0_0_296), .B2(
      n_0_0_108), .ZN(n_0_134));
   AOI22_X1 i_0_0_396 (.A1(n_0_0_85), .A2(n_0_37), .B1(n_0_0_86), .B2(
      read_data2[29]), .ZN(n_0_0_297));
   AOI22_X1 i_0_0_397 (.A1(n_0_0_88), .A2(n_0_67), .B1(n_0_0_89), .B2(
      read_data2[28]), .ZN(n_0_0_298));
   AND2_X1 i_0_0_398 (.A1(n_0_0_297), .A2(n_0_0_298), .ZN(n_0_0_299));
   INV_X1 i_0_0_399 (.A(n_0_0_173), .ZN(n_0_0_300));
   OAI22_X1 i_0_0_400 (.A1(n_0_0_299), .A2(shift[4]), .B1(n_0_0_300), .B2(
      n_0_0_69), .ZN(n_0_0_301));
   AOI22_X1 i_0_0_401 (.A1(n_0_0_301), .A2(n_0_0_142), .B1(n_0_0_235), .B2(
      shift[3]), .ZN(n_0_0_302));
   OAI22_X1 i_0_0_402 (.A1(n_0_0_302), .A2(shift[2]), .B1(n_0_0_268), .B2(
      n_0_0_70), .ZN(n_0_0_303));
   AOI22_X1 i_0_0_403 (.A1(n_0_0_303), .A2(n_0_0_101), .B1(n_0_0_287), .B2(
      shift[1]), .ZN(n_0_0_304));
   OAI22_X1 i_0_0_404 (.A1(n_0_0_304), .A2(n_0_0_108), .B1(n_0_0_296), .B2(
      n_0_0_109), .ZN(n_0_135));
   AOI22_X1 i_0_0_405 (.A1(n_0_0_85), .A2(n_0_38), .B1(n_0_0_88), .B2(n_0_68), 
      .ZN(n_0_0_305));
   AOI22_X1 i_0_0_406 (.A1(n_0_0_86), .A2(read_data2[30]), .B1(read_data2[29]), 
      .B2(n_0_0_89), .ZN(n_0_0_306));
   AND2_X1 i_0_0_407 (.A1(n_0_0_305), .A2(n_0_0_306), .ZN(n_0_0_307));
   INV_X1 i_0_0_408 (.A(n_0_0_179), .ZN(n_0_0_308));
   OAI22_X1 i_0_0_409 (.A1(n_0_0_307), .A2(shift[4]), .B1(n_0_0_308), .B2(
      n_0_0_69), .ZN(n_0_0_309));
   AOI22_X1 i_0_0_410 (.A1(n_0_0_309), .A2(n_0_0_142), .B1(n_0_0_242), .B2(
      shift[3]), .ZN(n_0_0_310));
   OAI22_X1 i_0_0_411 (.A1(n_0_0_277), .A2(n_0_0_70), .B1(n_0_0_310), .B2(
      shift[2]), .ZN(n_0_0_311));
   AOI22_X1 i_0_0_412 (.A1(n_0_0_311), .A2(n_0_0_101), .B1(n_0_0_295), .B2(
      shift[1]), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_413 (.A1(n_0_0_312), .A2(n_0_0_108), .B1(n_0_0_304), .B2(
      n_0_0_109), .ZN(n_0_136));
   AOI22_X1 i_0_0_414 (.A1(n_0_0_85), .A2(n_0_39), .B1(n_0_0_86), .B2(
      read_data2[31]), .ZN(n_0_0_313));
   INV_X1 i_0_0_415 (.A(n_0_0_313), .ZN(n_0_0_314));
   AOI221_X1 i_0_0_416 (.A(n_0_0_314), .B1(n_0_69), .B2(n_0_0_88), .C1(
      read_data2[30]), .C2(n_0_0_89), .ZN(n_0_0_315));
   INV_X1 i_0_0_417 (.A(n_0_0_185), .ZN(n_0_0_316));
   OAI22_X1 i_0_0_418 (.A1(n_0_0_315), .A2(shift[4]), .B1(n_0_0_316), .B2(
      n_0_0_69), .ZN(n_0_0_317));
   AOI22_X1 i_0_0_419 (.A1(n_0_0_317), .A2(n_0_0_142), .B1(shift[3]), .B2(
      n_0_0_249), .ZN(n_0_0_318));
   OAI22_X1 i_0_0_420 (.A1(n_0_0_318), .A2(shift[2]), .B1(n_0_0_286), .B2(
      n_0_0_70), .ZN(n_0_0_319));
   AOI22_X1 i_0_0_421 (.A1(n_0_0_319), .A2(n_0_0_101), .B1(n_0_0_303), .B2(
      shift[1]), .ZN(n_0_0_320));
   OAI22_X1 i_0_0_422 (.A1(n_0_0_320), .A2(n_0_0_108), .B1(n_0_0_312), .B2(
      n_0_0_109), .ZN(n_0_137));
   AOI221_X1 i_0_0_423 (.A(n_0_0_314), .B1(n_0_70), .B2(n_0_0_88), .C1(
      read_data2[31]), .C2(n_0_0_89), .ZN(n_0_0_321));
   NOR2_X1 i_0_0_424 (.A1(n_0_0_321), .A2(shift[4]), .ZN(n_0_0_322));
   INV_X1 i_0_0_425 (.A(n_0_0_322), .ZN(n_0_0_323));
   NOR2_X1 i_0_0_426 (.A1(n_0_0_323), .A2(shift[3]), .ZN(n_0_0_324));
   INV_X1 i_0_0_427 (.A(n_0_0_324), .ZN(n_0_0_325));
   NAND2_X1 i_0_0_428 (.A1(n_0_0_142), .A2(shift[4]), .ZN(n_0_0_326));
   OAI21_X1 i_0_0_429 (.A(n_0_0_325), .B1(n_0_0_192), .B2(n_0_0_326), .ZN(
      n_0_0_327));
   AOI21_X1 i_0_0_430 (.A(n_0_0_327), .B1(shift[3]), .B2(n_0_0_258), .ZN(
      n_0_0_328));
   OAI22_X1 i_0_0_431 (.A1(n_0_0_328), .A2(shift[2]), .B1(n_0_0_294), .B2(
      n_0_0_70), .ZN(n_0_0_329));
   AOI22_X1 i_0_0_432 (.A1(n_0_0_329), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_311), .ZN(n_0_0_330));
   OAI22_X1 i_0_0_433 (.A1(n_0_0_330), .A2(n_0_0_108), .B1(n_0_0_320), .B2(
      n_0_0_109), .ZN(n_0_138));
   NAND2_X1 i_0_0_434 (.A1(n_0_0_323), .A2(n_0_0_142), .ZN(n_0_0_331));
   NOR2_X1 i_0_0_435 (.A1(n_0_0_200), .A2(n_0_0_69), .ZN(n_0_0_332));
   OAI22_X1 i_0_0_436 (.A1(n_0_0_331), .A2(n_0_0_332), .B1(n_0_0_142), .B2(
      n_0_0_267), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_437 (.A1(n_0_0_333), .A2(shift[2]), .B1(n_0_0_70), .B2(
      n_0_0_302), .ZN(n_0_0_334));
   AOI22_X1 i_0_0_438 (.A1(n_0_0_334), .A2(n_0_0_101), .B1(n_0_0_319), .B2(
      shift[1]), .ZN(n_0_0_335));
   OAI22_X1 i_0_0_439 (.A1(n_0_0_330), .A2(n_0_0_109), .B1(n_0_0_335), .B2(
      n_0_0_108), .ZN(n_0_139));
   NOR2_X1 i_0_0_440 (.A1(n_0_0_211), .A2(n_0_0_69), .ZN(n_0_0_336));
   OAI22_X1 i_0_0_441 (.A1(n_0_0_331), .A2(n_0_0_336), .B1(n_0_0_142), .B2(
      n_0_0_276), .ZN(n_0_0_337));
   OAI22_X1 i_0_0_442 (.A1(n_0_0_337), .A2(shift[2]), .B1(n_0_0_310), .B2(
      n_0_0_70), .ZN(n_0_0_338));
   AOI22_X1 i_0_0_443 (.A1(n_0_0_329), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_338), .ZN(n_0_0_339));
   OAI22_X1 i_0_0_444 (.A1(n_0_0_339), .A2(n_0_0_108), .B1(n_0_0_335), .B2(
      n_0_0_109), .ZN(n_0_140));
   NOR2_X1 i_0_0_445 (.A1(n_0_0_219), .A2(n_0_0_69), .ZN(n_0_0_340));
   OAI22_X1 i_0_0_446 (.A1(n_0_0_331), .A2(n_0_0_340), .B1(n_0_0_142), .B2(
      n_0_0_285), .ZN(n_0_0_341));
   OAI22_X1 i_0_0_447 (.A1(n_0_0_341), .A2(shift[2]), .B1(n_0_0_318), .B2(
      n_0_0_70), .ZN(n_0_0_342));
   AOI22_X1 i_0_0_448 (.A1(n_0_0_101), .A2(n_0_0_342), .B1(n_0_0_334), .B2(
      shift[1]), .ZN(n_0_0_343));
   OAI22_X1 i_0_0_449 (.A1(n_0_0_339), .A2(n_0_0_109), .B1(n_0_0_343), .B2(
      n_0_0_108), .ZN(n_0_141));
   INV_X1 i_0_0_450 (.A(n_0_0_326), .ZN(n_0_0_344));
   AOI221_X1 i_0_0_451 (.A(n_0_0_324), .B1(n_0_0_226), .B2(n_0_0_344), .C1(
      shift[3]), .C2(n_0_0_293), .ZN(n_0_0_345));
   OAI22_X1 i_0_0_452 (.A1(n_0_0_345), .A2(shift[2]), .B1(n_0_0_328), .B2(
      n_0_0_70), .ZN(n_0_0_346));
   AOI22_X1 i_0_0_453 (.A1(n_0_0_346), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_338), .ZN(n_0_0_347));
   OAI22_X1 i_0_0_454 (.A1(n_0_0_347), .A2(n_0_0_108), .B1(n_0_0_343), .B2(
      n_0_0_109), .ZN(n_0_142));
   OAI21_X1 i_0_0_455 (.A(n_0_0_323), .B1(n_0_0_69), .B2(n_0_0_234), .ZN(
      n_0_0_348));
   OAI22_X1 i_0_0_456 (.A1(n_0_0_348), .A2(shift[3]), .B1(n_0_0_142), .B2(
      n_0_0_301), .ZN(n_0_0_349));
   AOI22_X1 i_0_0_457 (.A1(n_0_0_349), .A2(n_0_0_70), .B1(n_0_0_333), .B2(
      shift[2]), .ZN(n_0_0_350));
   AOI22_X1 i_0_0_458 (.A1(n_0_0_350), .A2(n_0_0_101), .B1(n_0_0_342), .B2(
      shift[1]), .ZN(n_0_0_351));
   OAI22_X1 i_0_0_459 (.A1(n_0_0_347), .A2(n_0_0_109), .B1(n_0_0_351), .B2(
      n_0_0_108), .ZN(n_0_143));
   OAI21_X1 i_0_0_460 (.A(n_0_0_323), .B1(n_0_0_69), .B2(n_0_0_241), .ZN(
      n_0_0_352));
   OAI22_X1 i_0_0_461 (.A1(n_0_0_352), .A2(shift[3]), .B1(n_0_0_142), .B2(
      n_0_0_309), .ZN(n_0_0_353));
   AOI22_X1 i_0_0_462 (.A1(n_0_0_353), .A2(n_0_0_70), .B1(n_0_0_337), .B2(
      shift[2]), .ZN(n_0_0_354));
   AOI22_X1 i_0_0_463 (.A1(n_0_0_346), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_354), .ZN(n_0_0_355));
   OAI22_X1 i_0_0_464 (.A1(n_0_0_355), .A2(n_0_0_108), .B1(n_0_0_351), .B2(
      n_0_0_109), .ZN(n_0_144));
   OAI21_X1 i_0_0_465 (.A(n_0_0_323), .B1(n_0_0_69), .B2(n_0_0_248), .ZN(
      n_0_0_356));
   OAI22_X1 i_0_0_466 (.A1(n_0_0_356), .A2(shift[3]), .B1(n_0_0_317), .B2(
      n_0_0_142), .ZN(n_0_0_357));
   AOI22_X1 i_0_0_467 (.A1(n_0_0_357), .A2(n_0_0_70), .B1(n_0_0_341), .B2(
      shift[2]), .ZN(n_0_0_358));
   OAI22_X1 i_0_0_468 (.A1(n_0_0_350), .A2(n_0_0_101), .B1(n_0_0_358), .B2(
      shift[1]), .ZN(n_0_0_359));
   OAI22_X1 i_0_0_469 (.A1(n_0_0_355), .A2(n_0_0_109), .B1(n_0_0_359), .B2(
      n_0_0_108), .ZN(n_0_145));
   OAI21_X1 i_0_0_470 (.A(n_0_0_323), .B1(n_0_0_256), .B2(n_0_0_326), .ZN(
      n_0_0_360));
   NAND2_X1 i_0_0_471 (.A1(shift[4]), .A2(shift[3]), .ZN(n_0_0_361));
   INV_X1 i_0_0_472 (.A(n_0_0_361), .ZN(n_0_0_362));
   AOI21_X1 i_0_0_473 (.A(n_0_0_360), .B1(n_0_0_191), .B2(n_0_0_362), .ZN(
      n_0_0_363));
   OAI22_X1 i_0_0_474 (.A1(n_0_0_345), .A2(n_0_0_70), .B1(shift[2]), .B2(
      n_0_0_363), .ZN(n_0_0_364));
   OAI22_X1 i_0_0_475 (.A1(n_0_0_364), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_354), .ZN(n_0_0_365));
   OAI22_X1 i_0_0_476 (.A1(n_0_0_365), .A2(n_0_0_108), .B1(n_0_0_359), .B2(
      n_0_0_109), .ZN(n_0_146));
   AOI221_X1 i_0_0_477 (.A(n_0_0_322), .B1(n_0_0_199), .B2(n_0_0_362), .C1(
      n_0_0_265), .C2(n_0_0_344), .ZN(n_0_0_366));
   AOI22_X1 i_0_0_478 (.A1(n_0_0_366), .A2(n_0_0_70), .B1(n_0_0_349), .B2(
      shift[2]), .ZN(n_0_0_367));
   OAI22_X1 i_0_0_479 (.A1(n_0_0_367), .A2(shift[1]), .B1(n_0_0_358), .B2(
      n_0_0_101), .ZN(n_0_0_368));
   OAI22_X1 i_0_0_480 (.A1(n_0_0_365), .A2(n_0_0_109), .B1(n_0_0_368), .B2(
      n_0_0_108), .ZN(n_0_147));
   AOI221_X1 i_0_0_481 (.A(n_0_0_322), .B1(n_0_0_210), .B2(n_0_0_362), .C1(
      n_0_0_274), .C2(n_0_0_344), .ZN(n_0_0_369));
   AOI22_X1 i_0_0_482 (.A1(n_0_0_369), .A2(n_0_0_70), .B1(n_0_0_353), .B2(
      shift[2]), .ZN(n_0_0_370));
   OAI22_X1 i_0_0_483 (.A1(n_0_0_364), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_370), .ZN(n_0_0_371));
   OAI22_X1 i_0_0_484 (.A1(n_0_0_371), .A2(n_0_0_108), .B1(n_0_0_368), .B2(
      n_0_0_109), .ZN(n_0_148));
   AOI221_X1 i_0_0_485 (.A(n_0_0_322), .B1(n_0_0_218), .B2(n_0_0_362), .C1(
      n_0_0_282), .C2(n_0_0_344), .ZN(n_0_0_372));
   AOI22_X1 i_0_0_486 (.A1(n_0_0_372), .A2(n_0_0_70), .B1(n_0_0_357), .B2(
      shift[2]), .ZN(n_0_0_373));
   OAI22_X1 i_0_0_487 (.A1(n_0_0_373), .A2(shift[1]), .B1(n_0_0_367), .B2(
      n_0_0_101), .ZN(n_0_0_374));
   OAI22_X1 i_0_0_488 (.A1(n_0_0_371), .A2(n_0_0_109), .B1(n_0_0_374), .B2(
      n_0_0_108), .ZN(n_0_149));
   OAI22_X1 i_0_0_489 (.A1(n_0_0_292), .A2(n_0_0_326), .B1(n_0_0_227), .B2(
      n_0_0_361), .ZN(n_0_0_375));
   NOR2_X1 i_0_0_490 (.A1(n_0_0_322), .A2(n_0_0_375), .ZN(n_0_0_376));
   OAI22_X1 i_0_0_491 (.A1(n_0_0_363), .A2(n_0_0_70), .B1(shift[2]), .B2(
      n_0_0_376), .ZN(n_0_0_377));
   OAI22_X1 i_0_0_492 (.A1(n_0_0_370), .A2(n_0_0_101), .B1(n_0_0_377), .B2(
      shift[1]), .ZN(n_0_0_378));
   OAI22_X1 i_0_0_493 (.A1(n_0_0_374), .A2(n_0_0_109), .B1(n_0_0_378), .B2(
      n_0_0_108), .ZN(n_0_150));
   OAI21_X1 i_0_0_494 (.A(n_0_0_323), .B1(n_0_0_69), .B2(n_0_0_299), .ZN(
      n_0_0_379));
   OAI22_X1 i_0_0_495 (.A1(n_0_0_348), .A2(n_0_0_142), .B1(n_0_0_379), .B2(
      shift[3]), .ZN(n_0_0_380));
   OAI22_X1 i_0_0_496 (.A1(shift[2]), .A2(n_0_0_380), .B1(n_0_0_366), .B2(
      n_0_0_70), .ZN(n_0_0_381));
   OAI22_X1 i_0_0_497 (.A1(n_0_0_381), .A2(shift[1]), .B1(n_0_0_373), .B2(
      n_0_0_101), .ZN(n_0_0_382));
   OAI22_X1 i_0_0_498 (.A1(n_0_0_382), .A2(n_0_0_108), .B1(n_0_0_378), .B2(
      n_0_0_109), .ZN(n_0_151));
   OAI21_X1 i_0_0_499 (.A(n_0_0_323), .B1(n_0_0_69), .B2(n_0_0_307), .ZN(
      n_0_0_383));
   OAI22_X1 i_0_0_500 (.A1(n_0_0_352), .A2(n_0_0_142), .B1(n_0_0_383), .B2(
      shift[3]), .ZN(n_0_0_384));
   OAI22_X1 i_0_0_501 (.A1(n_0_0_384), .A2(shift[2]), .B1(n_0_0_369), .B2(
      n_0_0_70), .ZN(n_0_0_385));
   AOI22_X1 i_0_0_502 (.A1(n_0_0_385), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_377), .ZN(n_0_0_386));
   OAI22_X1 i_0_0_503 (.A1(n_0_0_382), .A2(n_0_0_109), .B1(n_0_0_386), .B2(
      n_0_0_108), .ZN(n_0_152));
   NOR2_X1 i_0_0_504 (.A1(n_0_0_315), .A2(n_0_0_69), .ZN(n_0_0_387));
   OAI22_X1 i_0_0_505 (.A1(n_0_0_356), .A2(n_0_0_142), .B1(n_0_0_331), .B2(
      n_0_0_387), .ZN(n_0_0_388));
   OAI22_X1 i_0_0_506 (.A1(n_0_0_372), .A2(n_0_0_70), .B1(n_0_0_388), .B2(
      shift[2]), .ZN(n_0_0_389));
   AOI22_X1 i_0_0_507 (.A1(shift[1]), .A2(n_0_0_381), .B1(n_0_0_389), .B2(
      n_0_0_101), .ZN(n_0_0_390));
   OAI22_X1 i_0_0_508 (.A1(n_0_0_390), .A2(n_0_0_108), .B1(n_0_0_386), .B2(
      n_0_0_109), .ZN(n_0_153));
   NAND2_X1 i_0_0_509 (.A1(n_0_0_321), .A2(n_0_0_361), .ZN(n_0_0_391));
   OAI21_X1 i_0_0_510 (.A(n_0_0_391), .B1(n_0_0_255), .B2(n_0_0_361), .ZN(
      n_0_0_392));
   OAI22_X1 i_0_0_511 (.A1(n_0_0_376), .A2(n_0_0_70), .B1(n_0_0_392), .B2(
      shift[2]), .ZN(n_0_0_393));
   AOI22_X1 i_0_0_512 (.A1(n_0_0_385), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_393), .ZN(n_0_0_394));
   OAI22_X1 i_0_0_513 (.A1(n_0_0_390), .A2(n_0_0_109), .B1(n_0_0_394), .B2(
      n_0_0_108), .ZN(n_0_154));
   OAI21_X1 i_0_0_514 (.A(n_0_0_391), .B1(n_0_0_265), .B2(n_0_0_361), .ZN(
      n_0_0_395));
   AOI22_X1 i_0_0_515 (.A1(n_0_0_380), .A2(shift[2]), .B1(n_0_0_395), .B2(
      n_0_0_70), .ZN(n_0_0_396));
   AOI22_X1 i_0_0_516 (.A1(n_0_0_389), .A2(shift[1]), .B1(n_0_0_396), .B2(
      n_0_0_101), .ZN(n_0_0_397));
   OAI22_X1 i_0_0_517 (.A1(n_0_0_397), .A2(n_0_0_108), .B1(n_0_0_394), .B2(
      n_0_0_109), .ZN(n_0_155));
   OAI21_X1 i_0_0_518 (.A(n_0_0_391), .B1(n_0_0_274), .B2(n_0_0_361), .ZN(
      n_0_0_398));
   AOI22_X1 i_0_0_519 (.A1(n_0_0_384), .A2(shift[2]), .B1(n_0_0_70), .B2(
      n_0_0_398), .ZN(n_0_0_399));
   AOI22_X1 i_0_0_520 (.A1(n_0_0_399), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_393), .ZN(n_0_0_400));
   OAI22_X1 i_0_0_521 (.A1(n_0_0_397), .A2(n_0_0_109), .B1(n_0_0_400), .B2(
      n_0_0_108), .ZN(n_0_156));
   OAI211_X1 i_0_0_522 (.A(n_0_0_391), .B(n_0_0_70), .C1(n_0_0_282), .C2(
      n_0_0_361), .ZN(n_0_0_401));
   OAI21_X1 i_0_0_523 (.A(n_0_0_401), .B1(n_0_0_388), .B2(n_0_0_70), .ZN(
      n_0_0_402));
   OAI22_X1 i_0_0_524 (.A1(n_0_0_396), .A2(n_0_0_101), .B1(n_0_0_402), .B2(
      shift[1]), .ZN(n_0_0_403));
   OAI22_X1 i_0_0_525 (.A1(n_0_0_403), .A2(n_0_0_108), .B1(n_0_0_400), .B2(
      n_0_0_109), .ZN(n_0_157));
   NOR2_X1 i_0_0_526 (.A1(n_0_0_361), .A2(shift[2]), .ZN(n_0_0_404));
   INV_X1 i_0_0_527 (.A(n_0_0_404), .ZN(n_0_0_405));
   OAI22_X1 i_0_0_528 (.A1(n_0_0_392), .A2(n_0_0_404), .B1(n_0_0_292), .B2(
      n_0_0_405), .ZN(n_0_0_406));
   AOI22_X1 i_0_0_529 (.A1(n_0_0_399), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_406), .ZN(n_0_0_407));
   OAI22_X1 i_0_0_530 (.A1(n_0_0_403), .A2(n_0_0_109), .B1(n_0_0_407), .B2(
      n_0_0_108), .ZN(n_0_158));
   NAND2_X1 i_0_0_531 (.A1(n_0_0_379), .A2(shift[3]), .ZN(n_0_0_408));
   INV_X1 i_0_0_532 (.A(n_0_0_321), .ZN(n_0_0_409));
   AOI21_X1 i_0_0_533 (.A(shift[2]), .B1(n_0_0_409), .B2(n_0_0_142), .ZN(
      n_0_0_410));
   AOI22_X1 i_0_0_534 (.A1(n_0_0_408), .A2(n_0_0_410), .B1(shift[2]), .B2(
      n_0_0_395), .ZN(n_0_0_411));
   OAI22_X1 i_0_0_535 (.A1(n_0_0_402), .A2(n_0_0_101), .B1(n_0_0_411), .B2(
      shift[1]), .ZN(n_0_0_412));
   OAI22_X1 i_0_0_536 (.A1(n_0_0_407), .A2(n_0_0_109), .B1(n_0_0_412), .B2(
      n_0_0_108), .ZN(n_0_159));
   NAND2_X1 i_0_0_537 (.A1(n_0_0_383), .A2(shift[3]), .ZN(n_0_0_413));
   AOI22_X1 i_0_0_538 (.A1(n_0_0_413), .A2(n_0_0_410), .B1(shift[2]), .B2(
      n_0_0_398), .ZN(n_0_0_414));
   AOI22_X1 i_0_0_539 (.A1(n_0_0_414), .A2(n_0_0_101), .B1(shift[1]), .B2(
      n_0_0_406), .ZN(n_0_0_415));
   OAI22_X1 i_0_0_540 (.A1(n_0_0_412), .A2(n_0_0_109), .B1(n_0_0_415), .B2(
      n_0_0_108), .ZN(n_0_160));
   INV_X1 i_0_0_541 (.A(n_0_0_391), .ZN(n_0_0_416));
   NAND2_X1 i_0_0_542 (.A1(n_0_0_362), .A2(shift[2]), .ZN(n_0_0_417));
   INV_X1 i_0_0_543 (.A(n_0_0_417), .ZN(n_0_0_418));
   AOI221_X1 i_0_0_544 (.A(n_0_0_416), .B1(n_0_0_315), .B2(n_0_0_404), .C1(
      n_0_0_283), .C2(n_0_0_418), .ZN(n_0_0_419));
   OAI22_X1 i_0_0_545 (.A1(n_0_0_411), .A2(n_0_0_101), .B1(n_0_0_419), .B2(
      shift[1]), .ZN(n_0_0_420));
   OAI22_X1 i_0_0_546 (.A1(n_0_0_420), .A2(n_0_0_108), .B1(n_0_0_415), .B2(
      n_0_0_109), .ZN(n_0_161));
   NAND2_X1 i_0_0_547 (.A1(n_0_0_321), .A2(n_0_0_417), .ZN(n_0_0_421));
   INV_X1 i_0_0_548 (.A(n_0_0_421), .ZN(n_0_0_422));
   AOI21_X1 i_0_0_549 (.A(n_0_0_422), .B1(n_0_0_292), .B2(n_0_0_418), .ZN(
      n_0_0_423));
   AOI22_X1 i_0_0_550 (.A1(n_0_0_414), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_423), .ZN(n_0_0_424));
   OAI22_X1 i_0_0_551 (.A1(n_0_0_420), .A2(n_0_0_109), .B1(n_0_0_424), .B2(
      n_0_0_108), .ZN(n_0_162));
   NOR2_X1 i_0_0_552 (.A1(n_0_0_422), .A2(shift[1]), .ZN(n_0_0_425));
   INV_X1 i_0_0_553 (.A(n_0_0_425), .ZN(n_0_0_426));
   AOI21_X1 i_0_0_554 (.A(n_0_0_426), .B1(n_0_0_299), .B2(n_0_0_418), .ZN(
      n_0_0_427));
   AOI21_X1 i_0_0_555 (.A(n_0_0_427), .B1(n_0_0_419), .B2(shift[1]), .ZN(
      n_0_0_428));
   OAI22_X1 i_0_0_556 (.A1(n_0_0_428), .A2(n_0_0_108), .B1(n_0_0_424), .B2(
      n_0_0_109), .ZN(n_0_163));
   NAND2_X1 i_0_0_557 (.A1(n_0_0_307), .A2(n_0_0_418), .ZN(n_0_0_429));
   AOI22_X1 i_0_0_558 (.A1(n_0_0_423), .A2(shift[1]), .B1(n_0_0_425), .B2(
      n_0_0_429), .ZN(n_0_0_430));
   OAI22_X1 i_0_0_559 (.A1(n_0_0_428), .A2(n_0_0_109), .B1(n_0_0_430), .B2(
      n_0_0_108), .ZN(n_0_164));
   OAI22_X1 i_0_0_560 (.A1(n_0_0_315), .A2(shift[1]), .B1(n_0_0_101), .B2(
      n_0_0_299), .ZN(n_0_0_431));
   OAI21_X1 i_0_0_561 (.A(n_0_0_421), .B1(n_0_0_431), .B2(n_0_0_417), .ZN(
      n_0_0_432));
   OAI22_X1 i_0_0_562 (.A1(n_0_0_430), .A2(n_0_0_109), .B1(n_0_0_432), .B2(
      n_0_0_108), .ZN(n_0_165));
   NAND2_X1 i_0_0_563 (.A1(shift[2]), .A2(shift[1]), .ZN(n_0_0_433));
   INV_X1 i_0_0_564 (.A(n_0_0_433), .ZN(n_0_0_434));
   NAND2_X1 i_0_0_565 (.A1(n_0_0_434), .A2(shift[3]), .ZN(n_0_0_435));
   INV_X1 i_0_0_566 (.A(n_0_0_435), .ZN(n_0_0_436));
   NAND2_X1 i_0_0_567 (.A1(n_0_0_436), .A2(shift[4]), .ZN(n_0_0_437));
   NAND2_X1 i_0_0_568 (.A1(n_0_0_321), .A2(n_0_0_437), .ZN(n_0_0_438));
   OAI21_X1 i_0_0_569 (.A(n_0_0_438), .B1(n_0_0_101), .B2(n_0_0_429), .ZN(
      n_0_0_439));
   OAI22_X1 i_0_0_570 (.A1(n_0_0_432), .A2(n_0_0_109), .B1(n_0_0_439), .B2(
      n_0_0_108), .ZN(n_0_166));
   INV_X1 i_0_0_571 (.A(n_0_0_315), .ZN(n_0_0_440));
   OAI21_X1 i_0_0_572 (.A(n_0_0_438), .B1(n_0_0_440), .B2(n_0_0_437), .ZN(
      n_0_0_441));
   OAI22_X1 i_0_0_573 (.A1(n_0_0_439), .A2(n_0_0_109), .B1(n_0_0_441), .B2(
      n_0_0_108), .ZN(n_0_167));
   NOR2_X1 i_0_0_574 (.A1(n_0_0_321), .A2(n_0_0_94), .ZN(n_0_169));
   INV_X1 i_0_0_575 (.A(n_0_169), .ZN(n_0_0_442));
   AOI22_X1 i_0_0_576 (.A1(n_0_0_441), .A2(shift[0]), .B1(n_0_0_109), .B2(
      n_0_0_442), .ZN(n_0_168));
   OAI22_X1 i_0_0_577 (.A1(n_0_0_0), .A2(start_shift[0]), .B1(shift[0]), 
      .B2(start), .ZN(n_0_0_443));
   INV_X1 i_0_0_578 (.A(n_0_0_443), .ZN(n_0_170));
   INV_X1 i_0_0_579 (.A(start_shift[1]), .ZN(n_0_0_444));
   AOI22_X1 i_0_0_580 (.A1(n_0_0_444), .A2(start), .B1(n_0_0_0), .B2(shift[1]), 
      .ZN(n_0_171));
   OAI211_X1 i_0_0_581 (.A(n_0_0_433), .B(n_0_0_0), .C1(shift[2]), .C2(shift[1]), 
      .ZN(n_0_0_445));
   NAND2_X1 i_0_0_582 (.A1(start_shift[2]), .A2(start), .ZN(n_0_0_446));
   NAND2_X1 i_0_0_583 (.A1(n_0_0_445), .A2(n_0_0_446), .ZN(n_0_172));
   NAND2_X1 i_0_0_584 (.A1(start_shift[3]), .A2(start), .ZN(n_0_0_447));
   OAI21_X1 i_0_0_585 (.A(n_0_0_435), .B1(shift[3]), .B2(n_0_0_434), .ZN(
      n_0_0_448));
   OAI21_X1 i_0_0_586 (.A(n_0_0_447), .B1(n_0_0_448), .B2(start), .ZN(n_0_173));
   OAI211_X1 i_0_0_587 (.A(n_0_0_437), .B(n_0_0_0), .C1(shift[4]), .C2(n_0_0_436), 
      .ZN(n_0_0_449));
   NAND2_X1 i_0_0_588 (.A1(start), .A2(start_shift[4]), .ZN(n_0_0_450));
   NAND2_X1 i_0_0_589 (.A1(n_0_0_449), .A2(n_0_0_450), .ZN(n_0_174));
   DFF_X1 write_en_reg (.D(start), .CK(clk), .Q(write_en), .QN());
   DFF_X1 \c_reg[63]  (.D(n_0_125), .CK(clk), .Q(c[63]), .QN());
   DFF_X1 \c_reg[62]  (.D(n_0_124), .CK(clk), .Q(c[62]), .QN());
   DFF_X1 \c_reg[61]  (.D(n_0_123), .CK(clk), .Q(c[61]), .QN());
   DFF_X1 \c_reg[60]  (.D(n_0_122), .CK(clk), .Q(c[60]), .QN());
   DFF_X1 \c_reg[59]  (.D(n_0_121), .CK(clk), .Q(c[59]), .QN());
   DFF_X1 \c_reg[58]  (.D(n_0_120), .CK(clk), .Q(c[58]), .QN());
   DFF_X1 \c_reg[57]  (.D(n_0_119), .CK(clk), .Q(c[57]), .QN());
   DFF_X1 \c_reg[56]  (.D(n_0_118), .CK(clk), .Q(c[56]), .QN());
   DFF_X1 \c_reg[55]  (.D(n_0_117), .CK(clk), .Q(c[55]), .QN());
   DFF_X1 \c_reg[54]  (.D(n_0_116), .CK(clk), .Q(c[54]), .QN());
   DFF_X1 \c_reg[53]  (.D(n_0_115), .CK(clk), .Q(c[53]), .QN());
   DFF_X1 \c_reg[52]  (.D(n_0_114), .CK(clk), .Q(c[52]), .QN());
   DFF_X1 \c_reg[51]  (.D(n_0_113), .CK(clk), .Q(c[51]), .QN());
   DFF_X1 \c_reg[50]  (.D(n_0_112), .CK(clk), .Q(c[50]), .QN());
   DFF_X1 \c_reg[49]  (.D(n_0_111), .CK(clk), .Q(c[49]), .QN());
   DFF_X1 \c_reg[48]  (.D(n_0_110), .CK(clk), .Q(c[48]), .QN());
   DFF_X1 \c_reg[47]  (.D(n_0_109), .CK(clk), .Q(c[47]), .QN());
   DFF_X1 \c_reg[46]  (.D(n_0_108), .CK(clk), .Q(c[46]), .QN());
   DFF_X1 \c_reg[45]  (.D(n_0_107), .CK(clk), .Q(c[45]), .QN());
   DFF_X1 \c_reg[44]  (.D(n_0_106), .CK(clk), .Q(c[44]), .QN());
   DFF_X1 \c_reg[43]  (.D(n_0_105), .CK(clk), .Q(c[43]), .QN());
   DFF_X1 \c_reg[42]  (.D(n_0_104), .CK(clk), .Q(c[42]), .QN());
   DFF_X1 \c_reg[41]  (.D(n_0_103), .CK(clk), .Q(c[41]), .QN());
   DFF_X1 \c_reg[40]  (.D(n_0_102), .CK(clk), .Q(c[40]), .QN());
   DFF_X1 \c_reg[39]  (.D(n_0_101), .CK(clk), .Q(c[39]), .QN());
   DFF_X1 \c_reg[38]  (.D(n_0_100), .CK(clk), .Q(c[38]), .QN());
   DFF_X1 \c_reg[37]  (.D(n_0_99), .CK(clk), .Q(c[37]), .QN());
   DFF_X1 \c_reg[36]  (.D(n_0_98), .CK(clk), .Q(c[36]), .QN());
   DFF_X1 \c_reg[35]  (.D(n_0_97), .CK(clk), .Q(c[35]), .QN());
   DFF_X1 \c_reg[34]  (.D(n_0_96), .CK(clk), .Q(c[34]), .QN());
   DFF_X1 \c_reg[33]  (.D(n_0_95), .CK(clk), .Q(c[33]), .QN());
   DFF_X1 \c_reg[32]  (.D(n_0_94), .CK(clk), .Q(c[32]), .QN());
   DFF_X1 \c_reg[31]  (.D(n_0_93), .CK(clk), .Q(c[31]), .QN());
   DFF_X1 \c_reg[30]  (.D(n_0_92), .CK(clk), .Q(c[30]), .QN());
   DFF_X1 \c_reg[29]  (.D(n_0_91), .CK(clk), .Q(c[29]), .QN());
   DFF_X1 \c_reg[28]  (.D(n_0_90), .CK(clk), .Q(c[28]), .QN());
   DFF_X1 \c_reg[27]  (.D(n_0_89), .CK(clk), .Q(c[27]), .QN());
   DFF_X1 \c_reg[26]  (.D(n_0_88), .CK(clk), .Q(c[26]), .QN());
   DFF_X1 \c_reg[25]  (.D(n_0_87), .CK(clk), .Q(c[25]), .QN());
   DFF_X1 \c_reg[24]  (.D(n_0_86), .CK(clk), .Q(c[24]), .QN());
   DFF_X1 \c_reg[23]  (.D(n_0_85), .CK(clk), .Q(c[23]), .QN());
   DFF_X1 \c_reg[22]  (.D(n_0_84), .CK(clk), .Q(c[22]), .QN());
   DFF_X1 \c_reg[21]  (.D(n_0_83), .CK(clk), .Q(c[21]), .QN());
   DFF_X1 \c_reg[20]  (.D(n_0_82), .CK(clk), .Q(c[20]), .QN());
   DFF_X1 \c_reg[19]  (.D(n_0_81), .CK(clk), .Q(c[19]), .QN());
   DFF_X1 \c_reg[18]  (.D(n_0_80), .CK(clk), .Q(c[18]), .QN());
   DFF_X1 \c_reg[17]  (.D(n_0_79), .CK(clk), .Q(c[17]), .QN());
   DFF_X1 \c_reg[16]  (.D(n_0_78), .CK(clk), .Q(c[16]), .QN());
   DFF_X1 \c_reg[15]  (.D(n_0_77), .CK(clk), .Q(c[15]), .QN());
   DFF_X1 \c_reg[14]  (.D(n_0_76), .CK(clk), .Q(c[14]), .QN());
   DFF_X1 \c_reg[13]  (.D(n_0_75), .CK(clk), .Q(c[13]), .QN());
   DFF_X1 \c_reg[12]  (.D(n_0_74), .CK(clk), .Q(c[12]), .QN());
   DFF_X1 \c_reg[11]  (.D(n_0_73), .CK(clk), .Q(c[11]), .QN());
   DFF_X1 \c_reg[10]  (.D(n_0_72), .CK(clk), .Q(c[10]), .QN());
   DFF_X1 \c_reg[9]  (.D(n_0_71), .CK(clk), .Q(c[9]), .QN());
   DFF_X1 \c_reg[8]  (.D(n_0_8), .CK(clk), .Q(c[8]), .QN());
   DFF_X1 \c_reg[7]  (.D(n_0_7), .CK(clk), .Q(c[7]), .QN());
   DFF_X1 \c_reg[6]  (.D(n_0_6), .CK(clk), .Q(c[6]), .QN());
   DFF_X1 \c_reg[5]  (.D(n_0_5), .CK(clk), .Q(c[5]), .QN());
   DFF_X1 \c_reg[4]  (.D(n_0_4), .CK(clk), .Q(c[4]), .QN());
   DFF_X1 \c_reg[3]  (.D(n_0_3), .CK(clk), .Q(c[3]), .QN());
   DFF_X1 \c_reg[2]  (.D(n_0_2), .CK(clk), .Q(c[2]), .QN());
   DFF_X1 \c_reg[1]  (.D(n_0_1), .CK(clk), .Q(c[1]), .QN());
   DFF_X1 \c_reg[0]  (.D(n_0_0), .CK(clk), .Q(c[0]), .QN());
   DFF_X1 \shift_reg[4]  (.D(n_0_174), .CK(n_0_175), .Q(shift[4]), .QN());
   DFF_X1 \shift_reg[3]  (.D(n_0_173), .CK(n_0_175), .Q(shift[3]), .QN());
   DFF_X1 \shift_reg[2]  (.D(n_0_172), .CK(n_0_175), .Q(shift[2]), .QN());
   DFF_X1 \shift_reg[1]  (.D(n_0_171), .CK(n_0_175), .Q(shift[1]), .QN());
   DFF_X1 \shift_reg[0]  (.D(n_0_170), .CK(n_0_175), .Q(shift[0]), .QN());
   DFF_X1 \i_reg[4]  (.D(n_0_130), .CK(n_0_175), .Q(i[4]), .QN());
   DFF_X1 \i_reg[3]  (.D(n_0_129), .CK(n_0_175), .Q(i[3]), .QN());
   DFF_X1 \i_reg[2]  (.D(n_0_128), .CK(n_0_175), .Q(i[2]), .QN());
   DFF_X1 \i_reg[1]  (.D(n_0_127), .CK(n_0_175), .Q(i[1]), .QN());
   DFF_X1 \i_reg[0]  (.D(n_0_126), .CK(n_0_175), .Q(i[0]), .QN());
   CLKGATETST_X1 clk_gate_i_reg (.CK(clk), .E(n_0_131), .SE(1'b0), .GCK(n_0_175));
endmodule
