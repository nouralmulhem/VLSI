
// 	Wed Jan  4 14:44:47 2023
//	vlsi
//	localhost.localdomain

module datapath__0_142 (c, p_0, p_1);

output [63:0] p_1;
input [63:0] c;
input [63:0] p_0;
wire n_132;
wire n_200;
wire n_197;
wire n_0;
wire n_201;
wire n_198;
wire n_134;
wire n_130;
wire n_129;
wire n_127;
wire n_126;
wire n_124;
wire n_123;
wire n_121;
wire n_120;
wire n_118;
wire n_117;
wire n_115;
wire n_114;
wire n_112;
wire n_111;
wire n_109;
wire n_108;
wire n_106;
wire n_105;
wire n_103;
wire n_102;
wire n_100;
wire n_99;
wire n_97;
wire n_96;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_1;
wire n_202;
wire n_199;
wire n_137;
wire n_89;
wire n_88;
wire n_86;
wire n_85;
wire n_83;
wire n_82;
wire n_80;
wire n_79;
wire n_2;
wire n_139;
wire n_141;
wire n_78;
wire n_77;
wire n_3;
wire n_142;
wire n_143;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_4;
wire n_146;
wire n_148;
wire n_71;
wire n_70;
wire n_5;
wire n_149;
wire n_150;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_6;
wire n_153;
wire n_155;
wire n_64;
wire n_63;
wire n_7;
wire n_156;
wire n_157;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_8;
wire n_160;
wire n_162;
wire n_57;
wire n_56;
wire n_9;
wire n_163;
wire n_164;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_10;
wire n_167;
wire n_169;
wire n_50;
wire n_49;
wire n_11;
wire n_170;
wire n_171;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_12;
wire n_174;
wire n_176;
wire n_43;
wire n_42;
wire n_13;
wire n_177;
wire n_178;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_14;
wire n_181;
wire n_183;
wire n_36;
wire n_35;
wire n_15;
wire n_184;
wire n_185;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_16;
wire n_188;
wire n_190;
wire n_29;
wire n_28;
wire n_17;
wire n_191;
wire n_192;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_18;
wire n_194;
wire n_195;
wire n_21;
wire n_20;
wire n_19;
wire n_196;
wire n_22;
wire n_193;
wire n_27;
wire n_189;
wire n_187;
wire n_186;
wire n_34;
wire n_182;
wire n_180;
wire n_179;
wire n_41;
wire n_175;
wire n_173;
wire n_172;
wire n_48;
wire n_168;
wire n_166;
wire n_165;
wire n_55;
wire n_161;
wire n_159;
wire n_158;
wire n_62;
wire n_154;
wire n_152;
wire n_151;
wire n_69;
wire n_147;
wire n_145;
wire n_144;
wire n_76;
wire n_140;
wire n_138;
wire n_81;
wire n_84;
wire n_87;
wire n_136;
wire n_90;
wire n_135;
wire n_95;
wire n_98;
wire n_101;
wire n_104;
wire n_107;
wire n_110;
wire n_113;
wire n_116;
wire n_119;
wire n_122;
wire n_125;
wire n_128;
wire n_133;
wire n_131;


INV_X1 i_266 (.ZN (n_202), .A (c[16]));
INV_X1 i_265 (.ZN (n_201), .A (c[1]));
INV_X1 i_264 (.ZN (n_200), .A (c[0]));
INV_X1 i_263 (.ZN (n_199), .A (p_0[16]));
INV_X1 i_262 (.ZN (n_198), .A (p_0[1]));
INV_X1 i_261 (.ZN (n_197), .A (p_0[0]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (c[62]), .A2 (p_0[62]));
OAI21_X1 i_259 (.ZN (n_195), .A (n_196), .B1 (c[62]), .B2 (p_0[62]));
NAND2_X1 i_258 (.ZN (n_194), .A1 (c[61]), .A2 (p_0[61]));
NAND2_X1 i_257 (.ZN (n_193), .A1 (c[59]), .A2 (p_0[59]));
OAI21_X1 i_256 (.ZN (n_192), .A (n_193), .B1 (c[59]), .B2 (p_0[59]));
NAND2_X1 i_255 (.ZN (n_191), .A1 (c[58]), .A2 (p_0[58]));
XNOR2_X1 i_254 (.ZN (n_190), .A (c[57]), .B (p_0[57]));
INV_X1 i_253 (.ZN (n_189), .A (n_190));
NAND2_X1 i_252 (.ZN (n_188), .A1 (c[56]), .A2 (p_0[56]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (c[56]), .A2 (p_0[56]));
NAND2_X1 i_250 (.ZN (n_186), .A1 (c[54]), .A2 (p_0[54]));
OAI21_X1 i_249 (.ZN (n_185), .A (n_186), .B1 (c[54]), .B2 (p_0[54]));
NAND2_X1 i_248 (.ZN (n_184), .A1 (c[53]), .A2 (p_0[53]));
XNOR2_X1 i_247 (.ZN (n_183), .A (c[52]), .B (p_0[52]));
INV_X1 i_246 (.ZN (n_182), .A (n_183));
NAND2_X1 i_245 (.ZN (n_181), .A1 (c[51]), .A2 (p_0[51]));
NOR2_X1 i_244 (.ZN (n_180), .A1 (c[51]), .A2 (p_0[51]));
NAND2_X1 i_243 (.ZN (n_179), .A1 (c[49]), .A2 (p_0[49]));
OAI21_X1 i_242 (.ZN (n_178), .A (n_179), .B1 (c[49]), .B2 (p_0[49]));
NAND2_X1 i_241 (.ZN (n_177), .A1 (c[48]), .A2 (p_0[48]));
XNOR2_X1 i_240 (.ZN (n_176), .A (c[47]), .B (p_0[47]));
INV_X1 i_239 (.ZN (n_175), .A (n_176));
NAND2_X1 i_238 (.ZN (n_174), .A1 (c[46]), .A2 (p_0[46]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (c[46]), .A2 (p_0[46]));
NAND2_X1 i_236 (.ZN (n_172), .A1 (c[44]), .A2 (p_0[44]));
OAI21_X1 i_235 (.ZN (n_171), .A (n_172), .B1 (c[44]), .B2 (p_0[44]));
NAND2_X1 i_234 (.ZN (n_170), .A1 (c[43]), .A2 (p_0[43]));
XNOR2_X1 i_233 (.ZN (n_169), .A (c[42]), .B (p_0[42]));
INV_X1 i_232 (.ZN (n_168), .A (n_169));
NAND2_X1 i_231 (.ZN (n_167), .A1 (c[41]), .A2 (p_0[41]));
NOR2_X1 i_230 (.ZN (n_166), .A1 (c[41]), .A2 (p_0[41]));
NAND2_X1 i_229 (.ZN (n_165), .A1 (c[39]), .A2 (p_0[39]));
OAI21_X1 i_228 (.ZN (n_164), .A (n_165), .B1 (c[39]), .B2 (p_0[39]));
NAND2_X1 i_227 (.ZN (n_163), .A1 (c[38]), .A2 (p_0[38]));
XNOR2_X1 i_226 (.ZN (n_162), .A (c[37]), .B (p_0[37]));
INV_X1 i_225 (.ZN (n_161), .A (n_162));
NAND2_X1 i_224 (.ZN (n_160), .A1 (c[36]), .A2 (p_0[36]));
NOR2_X1 i_223 (.ZN (n_159), .A1 (c[36]), .A2 (p_0[36]));
NAND2_X1 i_222 (.ZN (n_158), .A1 (c[34]), .A2 (p_0[34]));
OAI21_X1 i_221 (.ZN (n_157), .A (n_158), .B1 (c[34]), .B2 (p_0[34]));
NAND2_X1 i_220 (.ZN (n_156), .A1 (c[33]), .A2 (p_0[33]));
XNOR2_X1 i_219 (.ZN (n_155), .A (c[32]), .B (p_0[32]));
INV_X1 i_218 (.ZN (n_154), .A (n_155));
NAND2_X1 i_217 (.ZN (n_153), .A1 (c[31]), .A2 (p_0[31]));
NOR2_X1 i_216 (.ZN (n_152), .A1 (c[31]), .A2 (p_0[31]));
NAND2_X1 i_215 (.ZN (n_151), .A1 (c[29]), .A2 (p_0[29]));
OAI21_X1 i_214 (.ZN (n_150), .A (n_151), .B1 (c[29]), .B2 (p_0[29]));
NAND2_X1 i_213 (.ZN (n_149), .A1 (c[28]), .A2 (p_0[28]));
XNOR2_X1 i_212 (.ZN (n_148), .A (c[27]), .B (p_0[27]));
INV_X1 i_211 (.ZN (n_147), .A (n_148));
NAND2_X1 i_210 (.ZN (n_146), .A1 (c[26]), .A2 (p_0[26]));
NOR2_X1 i_209 (.ZN (n_145), .A1 (c[26]), .A2 (p_0[26]));
NAND2_X1 i_208 (.ZN (n_144), .A1 (c[24]), .A2 (p_0[24]));
OAI21_X1 i_207 (.ZN (n_143), .A (n_144), .B1 (c[24]), .B2 (p_0[24]));
NAND2_X1 i_206 (.ZN (n_142), .A1 (c[23]), .A2 (p_0[23]));
XNOR2_X1 i_205 (.ZN (n_141), .A (c[22]), .B (p_0[22]));
INV_X1 i_204 (.ZN (n_140), .A (n_141));
NAND2_X1 i_203 (.ZN (n_139), .A1 (c[21]), .A2 (p_0[21]));
NOR2_X1 i_202 (.ZN (n_138), .A1 (c[21]), .A2 (p_0[21]));
XNOR2_X1 i_201 (.ZN (n_137), .A (c[17]), .B (p_0[17]));
INV_X1 i_200 (.ZN (n_136), .A (n_137));
NAND2_X1 i_199 (.ZN (n_135), .A1 (c[15]), .A2 (p_0[15]));
XNOR2_X1 i_198 (.ZN (n_134), .A (c[2]), .B (p_0[2]));
INV_X1 i_197 (.ZN (n_133), .A (n_134));
NOR2_X1 i_196 (.ZN (n_132), .A1 (n_200), .A2 (n_197));
AOI21_X1 i_195 (.ZN (n_131), .A (n_132), .B1 (c[1]), .B2 (p_0[1]));
AOI21_X1 i_194 (.ZN (n_130), .A (n_131), .B1 (n_201), .B2 (n_198));
AOI22_X1 i_193 (.ZN (n_129), .A1 (c[2]), .A2 (p_0[2]), .B1 (n_133), .B2 (n_130));
INV_X1 i_192 (.ZN (n_128), .A (n_129));
XOR2_X1 i_191 (.Z (n_127), .A (c[3]), .B (p_0[3]));
AOI22_X1 i_190 (.ZN (n_126), .A1 (c[3]), .A2 (p_0[3]), .B1 (n_128), .B2 (n_127));
INV_X1 i_189 (.ZN (n_125), .A (n_126));
XOR2_X1 i_188 (.Z (n_124), .A (c[4]), .B (p_0[4]));
AOI22_X1 i_187 (.ZN (n_123), .A1 (c[4]), .A2 (p_0[4]), .B1 (n_125), .B2 (n_124));
INV_X1 i_186 (.ZN (n_122), .A (n_123));
XOR2_X1 i_185 (.Z (n_121), .A (c[5]), .B (p_0[5]));
AOI22_X1 i_184 (.ZN (n_120), .A1 (c[5]), .A2 (p_0[5]), .B1 (n_122), .B2 (n_121));
INV_X1 i_183 (.ZN (n_119), .A (n_120));
XOR2_X1 i_182 (.Z (n_118), .A (c[6]), .B (p_0[6]));
AOI22_X2 i_181 (.ZN (n_117), .A1 (c[6]), .A2 (p_0[6]), .B1 (n_119), .B2 (n_118));
INV_X1 i_180 (.ZN (n_116), .A (n_117));
XOR2_X1 i_179 (.Z (n_115), .A (c[7]), .B (p_0[7]));
AOI22_X1 i_178 (.ZN (n_114), .A1 (c[7]), .A2 (p_0[7]), .B1 (n_116), .B2 (n_115));
INV_X1 i_177 (.ZN (n_113), .A (n_114));
XOR2_X1 i_176 (.Z (n_112), .A (c[8]), .B (p_0[8]));
AOI22_X1 i_175 (.ZN (n_111), .A1 (c[8]), .A2 (p_0[8]), .B1 (n_113), .B2 (n_112));
INV_X1 i_174 (.ZN (n_110), .A (n_111));
XOR2_X1 i_173 (.Z (n_109), .A (c[9]), .B (p_0[9]));
AOI22_X1 i_172 (.ZN (n_108), .A1 (c[9]), .A2 (p_0[9]), .B1 (n_110), .B2 (n_109));
INV_X1 i_171 (.ZN (n_107), .A (n_108));
XOR2_X1 i_170 (.Z (n_106), .A (c[10]), .B (p_0[10]));
AOI22_X1 i_169 (.ZN (n_105), .A1 (c[10]), .A2 (p_0[10]), .B1 (n_107), .B2 (n_106));
INV_X1 i_168 (.ZN (n_104), .A (n_105));
XOR2_X1 i_167 (.Z (n_103), .A (c[11]), .B (p_0[11]));
AOI22_X1 i_166 (.ZN (n_102), .A1 (c[11]), .A2 (p_0[11]), .B1 (n_104), .B2 (n_103));
INV_X1 i_165 (.ZN (n_101), .A (n_102));
XOR2_X1 i_164 (.Z (n_100), .A (c[12]), .B (p_0[12]));
AOI22_X2 i_163 (.ZN (n_99), .A1 (c[12]), .A2 (p_0[12]), .B1 (n_101), .B2 (n_100));
INV_X1 i_162 (.ZN (n_98), .A (n_99));
XOR2_X1 i_161 (.Z (n_97), .A (c[13]), .B (p_0[13]));
AOI22_X1 i_160 (.ZN (n_96), .A1 (c[13]), .A2 (p_0[13]), .B1 (n_98), .B2 (n_97));
INV_X1 i_159 (.ZN (n_95), .A (n_96));
XOR2_X1 i_158 (.Z (n_94), .A (c[14]), .B (p_0[14]));
AOI22_X1 i_157 (.ZN (n_93), .A1 (c[14]), .A2 (p_0[14]), .B1 (n_95), .B2 (n_94));
OAI21_X1 i_156 (.ZN (n_92), .A (n_135), .B1 (c[15]), .B2 (p_0[15]));
OAI21_X1 i_155 (.ZN (n_91), .A (n_135), .B1 (n_93), .B2 (n_92));
OAI21_X1 i_154 (.ZN (n_90), .A (n_91), .B1 (c[16]), .B2 (p_0[16]));
OAI21_X2 i_153 (.ZN (n_89), .A (n_90), .B1 (n_202), .B2 (n_199));
AOI22_X1 i_152 (.ZN (n_88), .A1 (c[17]), .A2 (p_0[17]), .B1 (n_136), .B2 (n_89));
INV_X1 i_151 (.ZN (n_87), .A (n_88));
XOR2_X1 i_150 (.Z (n_86), .A (c[18]), .B (p_0[18]));
AOI22_X1 i_149 (.ZN (n_85), .A1 (c[18]), .A2 (p_0[18]), .B1 (n_87), .B2 (n_86));
INV_X1 i_148 (.ZN (n_84), .A (n_85));
XOR2_X1 i_147 (.Z (n_83), .A (c[19]), .B (p_0[19]));
AOI22_X1 i_146 (.ZN (n_82), .A1 (c[19]), .A2 (p_0[19]), .B1 (n_84), .B2 (n_83));
INV_X1 i_145 (.ZN (n_81), .A (n_82));
XOR2_X1 i_144 (.Z (n_80), .A (c[20]), .B (p_0[20]));
AOI22_X1 i_143 (.ZN (n_79), .A1 (c[20]), .A2 (p_0[20]), .B1 (n_81), .B2 (n_80));
AOI21_X1 i_142 (.ZN (n_78), .A (n_138), .B1 (n_139), .B2 (n_79));
AOI22_X2 i_141 (.ZN (n_77), .A1 (c[22]), .A2 (p_0[22]), .B1 (n_140), .B2 (n_78));
NAND2_X1 i_140 (.ZN (n_76), .A1 (n_142), .A2 (n_77));
OAI21_X2 i_139 (.ZN (n_75), .A (n_76), .B1 (c[23]), .B2 (p_0[23]));
OAI21_X2 i_138 (.ZN (n_74), .A (n_144), .B1 (n_143), .B2 (n_75));
XOR2_X1 i_137 (.Z (n_73), .A (c[25]), .B (p_0[25]));
AOI22_X1 i_136 (.ZN (n_72), .A1 (c[25]), .A2 (p_0[25]), .B1 (n_74), .B2 (n_73));
AOI21_X2 i_135 (.ZN (n_71), .A (n_145), .B1 (n_146), .B2 (n_72));
AOI22_X1 i_134 (.ZN (n_70), .A1 (c[27]), .A2 (p_0[27]), .B1 (n_147), .B2 (n_71));
NAND2_X1 i_133 (.ZN (n_69), .A1 (n_149), .A2 (n_70));
OAI21_X2 i_132 (.ZN (n_68), .A (n_69), .B1 (c[28]), .B2 (p_0[28]));
OAI21_X2 i_131 (.ZN (n_67), .A (n_151), .B1 (n_150), .B2 (n_68));
XOR2_X1 i_130 (.Z (n_66), .A (c[30]), .B (p_0[30]));
AOI22_X2 i_129 (.ZN (n_65), .A1 (c[30]), .A2 (p_0[30]), .B1 (n_67), .B2 (n_66));
AOI21_X2 i_128 (.ZN (n_64), .A (n_152), .B1 (n_153), .B2 (n_65));
AOI22_X1 i_127 (.ZN (n_63), .A1 (c[32]), .A2 (p_0[32]), .B1 (n_154), .B2 (n_64));
NAND2_X1 i_126 (.ZN (n_62), .A1 (n_156), .A2 (n_63));
OAI21_X2 i_125 (.ZN (n_61), .A (n_62), .B1 (c[33]), .B2 (p_0[33]));
OAI21_X2 i_124 (.ZN (n_60), .A (n_158), .B1 (n_157), .B2 (n_61));
XOR2_X1 i_123 (.Z (n_59), .A (c[35]), .B (p_0[35]));
AOI22_X1 i_122 (.ZN (n_58), .A1 (c[35]), .A2 (p_0[35]), .B1 (n_60), .B2 (n_59));
AOI21_X2 i_121 (.ZN (n_57), .A (n_159), .B1 (n_160), .B2 (n_58));
AOI22_X1 i_120 (.ZN (n_56), .A1 (c[37]), .A2 (p_0[37]), .B1 (n_161), .B2 (n_57));
NAND2_X1 i_119 (.ZN (n_55), .A1 (n_163), .A2 (n_56));
OAI21_X2 i_118 (.ZN (n_54), .A (n_55), .B1 (c[38]), .B2 (p_0[38]));
OAI21_X2 i_117 (.ZN (n_53), .A (n_165), .B1 (n_164), .B2 (n_54));
XOR2_X1 i_116 (.Z (n_52), .A (c[40]), .B (p_0[40]));
AOI22_X1 i_115 (.ZN (n_51), .A1 (c[40]), .A2 (p_0[40]), .B1 (n_53), .B2 (n_52));
AOI21_X2 i_114 (.ZN (n_50), .A (n_166), .B1 (n_167), .B2 (n_51));
AOI22_X1 i_113 (.ZN (n_49), .A1 (c[42]), .A2 (p_0[42]), .B1 (n_168), .B2 (n_50));
NAND2_X1 i_112 (.ZN (n_48), .A1 (n_170), .A2 (n_49));
OAI21_X2 i_111 (.ZN (n_47), .A (n_48), .B1 (c[43]), .B2 (p_0[43]));
OAI21_X1 i_110 (.ZN (n_46), .A (n_172), .B1 (n_171), .B2 (n_47));
XOR2_X1 i_109 (.Z (n_45), .A (c[45]), .B (p_0[45]));
AOI22_X1 i_108 (.ZN (n_44), .A1 (c[45]), .A2 (p_0[45]), .B1 (n_46), .B2 (n_45));
AOI21_X2 i_107 (.ZN (n_43), .A (n_173), .B1 (n_174), .B2 (n_44));
AOI22_X1 i_106 (.ZN (n_42), .A1 (c[47]), .A2 (p_0[47]), .B1 (n_175), .B2 (n_43));
NAND2_X1 i_105 (.ZN (n_41), .A1 (n_177), .A2 (n_42));
OAI21_X1 i_104 (.ZN (n_40), .A (n_41), .B1 (c[48]), .B2 (p_0[48]));
OAI21_X1 i_103 (.ZN (n_39), .A (n_179), .B1 (n_178), .B2 (n_40));
XOR2_X1 i_102 (.Z (n_38), .A (c[50]), .B (p_0[50]));
AOI22_X1 i_101 (.ZN (n_37), .A1 (c[50]), .A2 (p_0[50]), .B1 (n_39), .B2 (n_38));
AOI21_X1 i_100 (.ZN (n_36), .A (n_180), .B1 (n_181), .B2 (n_37));
AOI22_X1 i_99 (.ZN (n_35), .A1 (c[52]), .A2 (p_0[52]), .B1 (n_182), .B2 (n_36));
NAND2_X1 i_98 (.ZN (n_34), .A1 (n_184), .A2 (n_35));
OAI21_X1 i_97 (.ZN (n_33), .A (n_34), .B1 (c[53]), .B2 (p_0[53]));
OAI21_X1 i_96 (.ZN (n_32), .A (n_186), .B1 (n_185), .B2 (n_33));
XOR2_X1 i_95 (.Z (n_31), .A (c[55]), .B (p_0[55]));
AOI22_X1 i_94 (.ZN (n_30), .A1 (c[55]), .A2 (p_0[55]), .B1 (n_32), .B2 (n_31));
AOI21_X1 i_93 (.ZN (n_29), .A (n_187), .B1 (n_188), .B2 (n_30));
AOI22_X1 i_92 (.ZN (n_28), .A1 (c[57]), .A2 (p_0[57]), .B1 (n_189), .B2 (n_29));
NAND2_X1 i_91 (.ZN (n_27), .A1 (n_191), .A2 (n_28));
OAI21_X1 i_90 (.ZN (n_26), .A (n_27), .B1 (c[58]), .B2 (p_0[58]));
OAI21_X1 i_89 (.ZN (n_25), .A (n_193), .B1 (n_192), .B2 (n_26));
XOR2_X1 i_88 (.Z (n_24), .A (c[60]), .B (p_0[60]));
AOI22_X1 i_87 (.ZN (n_23), .A1 (c[60]), .A2 (p_0[60]), .B1 (n_25), .B2 (n_24));
NAND2_X1 i_86 (.ZN (n_22), .A1 (n_194), .A2 (n_23));
OAI21_X1 i_85 (.ZN (n_21), .A (n_22), .B1 (c[61]), .B2 (p_0[61]));
OAI21_X1 i_84 (.ZN (n_20), .A (n_196), .B1 (n_195), .B2 (n_21));
XOR2_X1 i_83 (.Z (n_19), .A (c[63]), .B (p_0[63]));
XOR2_X1 i_82 (.Z (p_1[63]), .A (n_20), .B (n_19));
XOR2_X1 i_81 (.Z (p_1[62]), .A (n_195), .B (n_21));
OAI21_X1 i_80 (.ZN (n_18), .A (n_194), .B1 (c[61]), .B2 (p_0[61]));
XOR2_X1 i_79 (.Z (p_1[61]), .A (n_23), .B (n_18));
XOR2_X1 i_78 (.Z (p_1[60]), .A (n_25), .B (n_24));
XOR2_X1 i_77 (.Z (p_1[59]), .A (n_192), .B (n_26));
OAI21_X1 i_76 (.ZN (n_17), .A (n_191), .B1 (c[58]), .B2 (p_0[58]));
XOR2_X1 i_75 (.Z (p_1[58]), .A (n_28), .B (n_17));
XNOR2_X1 i_74 (.ZN (p_1[57]), .A (n_190), .B (n_29));
OAI21_X1 i_73 (.ZN (n_16), .A (n_188), .B1 (c[56]), .B2 (p_0[56]));
XOR2_X1 i_72 (.Z (p_1[56]), .A (n_30), .B (n_16));
XOR2_X1 i_71 (.Z (p_1[55]), .A (n_32), .B (n_31));
XOR2_X1 i_70 (.Z (p_1[54]), .A (n_185), .B (n_33));
OAI21_X1 i_69 (.ZN (n_15), .A (n_184), .B1 (c[53]), .B2 (p_0[53]));
XOR2_X1 i_68 (.Z (p_1[53]), .A (n_35), .B (n_15));
XNOR2_X1 i_67 (.ZN (p_1[52]), .A (n_183), .B (n_36));
OAI21_X1 i_66 (.ZN (n_14), .A (n_181), .B1 (c[51]), .B2 (p_0[51]));
XOR2_X1 i_65 (.Z (p_1[51]), .A (n_37), .B (n_14));
XOR2_X1 i_64 (.Z (p_1[50]), .A (n_39), .B (n_38));
XOR2_X1 i_63 (.Z (p_1[49]), .A (n_178), .B (n_40));
OAI21_X1 i_62 (.ZN (n_13), .A (n_177), .B1 (c[48]), .B2 (p_0[48]));
XOR2_X1 i_61 (.Z (p_1[48]), .A (n_42), .B (n_13));
XNOR2_X1 i_60 (.ZN (p_1[47]), .A (n_176), .B (n_43));
OAI21_X1 i_59 (.ZN (n_12), .A (n_174), .B1 (c[46]), .B2 (p_0[46]));
XOR2_X1 i_58 (.Z (p_1[46]), .A (n_44), .B (n_12));
XOR2_X1 i_57 (.Z (p_1[45]), .A (n_46), .B (n_45));
XOR2_X1 i_56 (.Z (p_1[44]), .A (n_171), .B (n_47));
OAI21_X1 i_55 (.ZN (n_11), .A (n_170), .B1 (c[43]), .B2 (p_0[43]));
XOR2_X1 i_54 (.Z (p_1[43]), .A (n_49), .B (n_11));
XNOR2_X1 i_53 (.ZN (p_1[42]), .A (n_169), .B (n_50));
OAI21_X1 i_52 (.ZN (n_10), .A (n_167), .B1 (c[41]), .B2 (p_0[41]));
XOR2_X1 i_51 (.Z (p_1[41]), .A (n_51), .B (n_10));
XOR2_X1 i_50 (.Z (p_1[40]), .A (n_53), .B (n_52));
XOR2_X1 i_49 (.Z (p_1[39]), .A (n_164), .B (n_54));
OAI21_X1 i_48 (.ZN (n_9), .A (n_163), .B1 (c[38]), .B2 (p_0[38]));
XOR2_X1 i_47 (.Z (p_1[38]), .A (n_56), .B (n_9));
XNOR2_X1 i_46 (.ZN (p_1[37]), .A (n_162), .B (n_57));
OAI21_X1 i_45 (.ZN (n_8), .A (n_160), .B1 (c[36]), .B2 (p_0[36]));
XOR2_X1 i_44 (.Z (p_1[36]), .A (n_58), .B (n_8));
XOR2_X1 i_43 (.Z (p_1[35]), .A (n_60), .B (n_59));
XOR2_X1 i_42 (.Z (p_1[34]), .A (n_157), .B (n_61));
OAI21_X1 i_41 (.ZN (n_7), .A (n_156), .B1 (c[33]), .B2 (p_0[33]));
XOR2_X1 i_40 (.Z (p_1[33]), .A (n_63), .B (n_7));
XNOR2_X1 i_39 (.ZN (p_1[32]), .A (n_155), .B (n_64));
OAI21_X1 i_38 (.ZN (n_6), .A (n_153), .B1 (c[31]), .B2 (p_0[31]));
XOR2_X1 i_37 (.Z (p_1[31]), .A (n_65), .B (n_6));
XOR2_X1 i_36 (.Z (p_1[30]), .A (n_67), .B (n_66));
XOR2_X1 i_35 (.Z (p_1[29]), .A (n_150), .B (n_68));
OAI21_X1 i_34 (.ZN (n_5), .A (n_149), .B1 (c[28]), .B2 (p_0[28]));
XOR2_X1 i_33 (.Z (p_1[28]), .A (n_70), .B (n_5));
XNOR2_X1 i_32 (.ZN (p_1[27]), .A (n_148), .B (n_71));
OAI21_X1 i_31 (.ZN (n_4), .A (n_146), .B1 (c[26]), .B2 (p_0[26]));
XOR2_X1 i_30 (.Z (p_1[26]), .A (n_72), .B (n_4));
XOR2_X1 i_29 (.Z (p_1[25]), .A (n_74), .B (n_73));
XOR2_X1 i_28 (.Z (p_1[24]), .A (n_143), .B (n_75));
OAI21_X1 i_27 (.ZN (n_3), .A (n_142), .B1 (c[23]), .B2 (p_0[23]));
XOR2_X1 i_26 (.Z (p_1[23]), .A (n_77), .B (n_3));
XNOR2_X1 i_25 (.ZN (p_1[22]), .A (n_141), .B (n_78));
OAI21_X1 i_24 (.ZN (n_2), .A (n_139), .B1 (c[21]), .B2 (p_0[21]));
XOR2_X1 i_23 (.Z (p_1[21]), .A (n_79), .B (n_2));
XNOR2_X1 i_22 (.ZN (p_1[20]), .A (n_82), .B (n_80));
XNOR2_X1 i_21 (.ZN (p_1[19]), .A (n_85), .B (n_83));
XNOR2_X1 i_20 (.ZN (p_1[18]), .A (n_88), .B (n_86));
XNOR2_X1 i_19 (.ZN (p_1[17]), .A (n_137), .B (n_89));
OAI22_X1 i_18 (.ZN (n_1), .A1 (c[16]), .A2 (p_0[16]), .B1 (n_202), .B2 (n_199));
XNOR2_X1 i_17 (.ZN (p_1[16]), .A (n_91), .B (n_1));
XOR2_X1 i_16 (.Z (p_1[15]), .A (n_93), .B (n_92));
XNOR2_X1 i_15 (.ZN (p_1[14]), .A (n_96), .B (n_94));
XNOR2_X1 i_14 (.ZN (p_1[13]), .A (n_99), .B (n_97));
XNOR2_X1 i_13 (.ZN (p_1[12]), .A (n_102), .B (n_100));
XNOR2_X1 i_12 (.ZN (p_1[11]), .A (n_105), .B (n_103));
XNOR2_X1 i_11 (.ZN (p_1[10]), .A (n_108), .B (n_106));
XNOR2_X1 i_10 (.ZN (p_1[9]), .A (n_111), .B (n_109));
XNOR2_X1 i_9 (.ZN (p_1[8]), .A (n_114), .B (n_112));
XNOR2_X1 i_8 (.ZN (p_1[7]), .A (n_117), .B (n_115));
XNOR2_X1 i_7 (.ZN (p_1[6]), .A (n_120), .B (n_118));
XNOR2_X1 i_6 (.ZN (p_1[5]), .A (n_123), .B (n_121));
XNOR2_X1 i_5 (.ZN (p_1[4]), .A (n_126), .B (n_124));
XNOR2_X1 i_4 (.ZN (p_1[3]), .A (n_129), .B (n_127));
XNOR2_X1 i_3 (.ZN (p_1[2]), .A (n_134), .B (n_130));
OAI22_X1 i_2 (.ZN (n_0), .A1 (n_201), .A2 (n_198), .B1 (c[1]), .B2 (p_0[1]));
XNOR2_X1 i_1 (.ZN (p_1[1]), .A (n_132), .B (n_0));
AOI21_X1 i_0 (.ZN (p_1[0]), .A (n_132), .B1 (n_200), .B2 (n_197));

endmodule //datapath__0_142

module datapath__0_128 (p_0, p_1);

output [32:0] p_0;
input [32:0] p_1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (p_1[25]));
INV_X1 i_63 (.ZN (n_32), .A (p_1[21]));
INV_X1 i_62 (.ZN (n_31), .A (p_1[14]));
INV_X1 i_61 (.ZN (n_30), .A (p_1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (p_1[2]), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (p_1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (p_1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (p_1[5]), .A3 (p_1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (p_1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (p_1[8]), .A3 (p_1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (p_1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (p_1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (p_1[12]), .A3 (p_1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (p_1[15]), .A3 (p_1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (p_1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (p_1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]), .A4 (p_1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (p_1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (p_1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (p_1[23]), .A3 (p_1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (p_1[26]), .A3 (p_1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (p_1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]), .A4 (p_1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (p_1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (p_1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (p_1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (p_1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (p_1[27]), .B1 (n_9), .B2 (p_1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (p_1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (p_1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (p_1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (p_1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (p_1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (p_1[16]), .B1 (n_19), .B2 (p_1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (p_1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (p_1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (p_1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (p_1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (p_1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (p_1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[9]), .B1 (n_25), .B2 (p_1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (p_1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (p_1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[6]), .B1 (n_27), .B2 (p_1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (p_1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (p_1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (p_1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[2]), .B1 (p_1[1]), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (p_1[1]), .B (p_1[0]));

endmodule //datapath__0_128

module datapath (p_0, read_data2);

output [31:0] p_0;
input [31:0] read_data2;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (read_data2[25]));
INV_X1 i_63 (.ZN (n_32), .A (read_data2[21]));
INV_X1 i_62 (.ZN (n_31), .A (read_data2[14]));
INV_X1 i_61 (.ZN (n_30), .A (read_data2[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (read_data2[2]), .A2 (read_data2[1]), .A3 (read_data2[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (read_data2[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (read_data2[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (read_data2[5]), .A3 (read_data2[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (read_data2[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (read_data2[8]), .A3 (read_data2[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (read_data2[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (read_data2[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (read_data2[12]), .A3 (read_data2[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (read_data2[15]), .A3 (read_data2[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (read_data2[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (read_data2[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (read_data2[18]), .A3 (read_data2[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (read_data2[18]), .A3 (read_data2[19]), .A4 (read_data2[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (read_data2[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (read_data2[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (read_data2[23]), .A3 (read_data2[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (read_data2[26]), .A3 (read_data2[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (read_data2[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (read_data2[28]), .A3 (read_data2[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (read_data2[28]), .A3 (read_data2[29]), .A4 (read_data2[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (read_data2[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (read_data2[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (read_data2[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (read_data2[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (read_data2[27]), .B1 (n_9), .B2 (read_data2[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (read_data2[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (read_data2[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (read_data2[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (read_data2[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (read_data2[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (read_data2[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (read_data2[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (read_data2[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (read_data2[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (read_data2[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (read_data2[16]), .B1 (n_19), .B2 (read_data2[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (read_data2[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (read_data2[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (read_data2[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (read_data2[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (read_data2[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (read_data2[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (read_data2[9]), .B1 (n_25), .B2 (read_data2[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (read_data2[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (read_data2[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (read_data2[6]), .B1 (n_27), .B2 (read_data2[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (read_data2[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (read_data2[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (read_data2[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (read_data2[2]), .B1 (read_data2[1]), .B2 (read_data2[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (read_data2[1]), .B (read_data2[0]));

endmodule //datapath

module regFile64 (clk__CTS_1_PP_0, read_data, write_en, write_data, clk);

output [63:0] read_data;
input clk;
input [63:0] write_data;
input write_en;
input clk__CTS_1_PP_0;
wire CTS_n_tid1_8;
wire CTS_n_tid1_7;


DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid1_7), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid1_7), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid1_7), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid1_7), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid1_7), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid1_7), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid1_7), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid1_7), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid1_7), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid1_7), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid1_7), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid1_7), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid1_7), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid1_7), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid1_7), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid1_7), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid1_7), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid1_7), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid1_7), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid1_7), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid1_7), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid1_7), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid1_7), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid1_7), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid1_7), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid1_7), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid1_7), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid1_7), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid1_7), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid1_7), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid1_7), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid1_7), .D (write_data[31]));
DFF_X1 \my_reg_reg[32]  (.Q (read_data[32]), .CK (CTS_n_tid1_7), .D (write_data[32]));
DFF_X1 \my_reg_reg[33]  (.Q (read_data[33]), .CK (CTS_n_tid1_7), .D (write_data[33]));
DFF_X1 \my_reg_reg[34]  (.Q (read_data[34]), .CK (CTS_n_tid1_7), .D (write_data[34]));
DFF_X1 \my_reg_reg[35]  (.Q (read_data[35]), .CK (CTS_n_tid1_7), .D (write_data[35]));
DFF_X1 \my_reg_reg[36]  (.Q (read_data[36]), .CK (CTS_n_tid1_7), .D (write_data[36]));
DFF_X1 \my_reg_reg[37]  (.Q (read_data[37]), .CK (CTS_n_tid1_7), .D (write_data[37]));
DFF_X1 \my_reg_reg[38]  (.Q (read_data[38]), .CK (CTS_n_tid1_7), .D (write_data[38]));
DFF_X1 \my_reg_reg[39]  (.Q (read_data[39]), .CK (CTS_n_tid1_7), .D (write_data[39]));
DFF_X1 \my_reg_reg[40]  (.Q (read_data[40]), .CK (CTS_n_tid1_7), .D (write_data[40]));
DFF_X1 \my_reg_reg[41]  (.Q (read_data[41]), .CK (CTS_n_tid1_7), .D (write_data[41]));
DFF_X1 \my_reg_reg[42]  (.Q (read_data[42]), .CK (CTS_n_tid1_7), .D (write_data[42]));
DFF_X1 \my_reg_reg[43]  (.Q (read_data[43]), .CK (CTS_n_tid1_7), .D (write_data[43]));
DFF_X1 \my_reg_reg[44]  (.Q (read_data[44]), .CK (CTS_n_tid1_7), .D (write_data[44]));
DFF_X1 \my_reg_reg[45]  (.Q (read_data[45]), .CK (CTS_n_tid1_7), .D (write_data[45]));
DFF_X1 \my_reg_reg[46]  (.Q (read_data[46]), .CK (CTS_n_tid1_7), .D (write_data[46]));
DFF_X1 \my_reg_reg[47]  (.Q (read_data[47]), .CK (CTS_n_tid1_7), .D (write_data[47]));
DFF_X1 \my_reg_reg[48]  (.Q (read_data[48]), .CK (CTS_n_tid1_7), .D (write_data[48]));
DFF_X1 \my_reg_reg[49]  (.Q (read_data[49]), .CK (CTS_n_tid1_7), .D (write_data[49]));
DFF_X1 \my_reg_reg[50]  (.Q (read_data[50]), .CK (CTS_n_tid1_7), .D (write_data[50]));
DFF_X1 \my_reg_reg[51]  (.Q (read_data[51]), .CK (CTS_n_tid1_7), .D (write_data[51]));
DFF_X1 \my_reg_reg[52]  (.Q (read_data[52]), .CK (CTS_n_tid1_7), .D (write_data[52]));
DFF_X1 \my_reg_reg[53]  (.Q (read_data[53]), .CK (CTS_n_tid1_7), .D (write_data[53]));
DFF_X1 \my_reg_reg[54]  (.Q (read_data[54]), .CK (CTS_n_tid1_7), .D (write_data[54]));
DFF_X1 \my_reg_reg[55]  (.Q (read_data[55]), .CK (CTS_n_tid1_7), .D (write_data[55]));
DFF_X1 \my_reg_reg[56]  (.Q (read_data[56]), .CK (CTS_n_tid1_7), .D (write_data[56]));
DFF_X1 \my_reg_reg[57]  (.Q (read_data[57]), .CK (CTS_n_tid1_7), .D (write_data[57]));
DFF_X1 \my_reg_reg[58]  (.Q (read_data[58]), .CK (CTS_n_tid1_7), .D (write_data[58]));
DFF_X1 \my_reg_reg[59]  (.Q (read_data[59]), .CK (CTS_n_tid1_7), .D (write_data[59]));
DFF_X1 \my_reg_reg[60]  (.Q (read_data[60]), .CK (CTS_n_tid1_7), .D (write_data[60]));
DFF_X1 \my_reg_reg[61]  (.Q (read_data[61]), .CK (CTS_n_tid1_7), .D (write_data[61]));
DFF_X1 \my_reg_reg[62]  (.Q (read_data[62]), .CK (CTS_n_tid1_7), .D (write_data[62]));
CLKBUF_X3 CTS_L4_c_tid1_4 (.Z (CTS_n_tid1_7), .A (CTS_n_tid1_8));
DFF_X1 \my_reg_reg[63]  (.Q (read_data[63]), .CK (CTS_n_tid1_7), .D (write_data[63]));
INV_X4 CTS_L3_c_tid1_5 (.ZN (CTS_n_tid1_8), .A (clk__CTS_1_PP_0));

endmodule //regFile64

module regFile (clk__CTS_1_PP_0, clk__CTS_1_PP_3, clk__CTS_1_PP_4, read_data, read_data2, 
    write_en, write_data, write_data2, clk);

output [31:0] read_data2;
output [31:0] read_data;
output clk__CTS_1_PP_0;
output clk__CTS_1_PP_3;
input clk;
input [31:0] write_data2;
input [31:0] write_data;
input write_en;
input clk__CTS_1_PP_4;
wire CTS_n_tid1_5;
wire CTS_n_tid1_6;


CLKGATETST_X8 clk_gate_my_reg_reg (.GCK (CTS_n_tid1_6), .CK (clk__CTS_1_PP_0), .E (write_en), .SE (1'b0 ));
DFF_X1 \my_reg_reg[0]  (.Q (read_data[0]), .CK (CTS_n_tid1_5), .D (write_data[0]));
DFF_X1 \my_reg_reg[1]  (.Q (read_data[1]), .CK (CTS_n_tid1_5), .D (write_data[1]));
DFF_X1 \my_reg_reg[2]  (.Q (read_data[2]), .CK (CTS_n_tid1_5), .D (write_data[2]));
DFF_X1 \my_reg_reg[3]  (.Q (read_data[3]), .CK (CTS_n_tid1_5), .D (write_data[3]));
DFF_X1 \my_reg_reg[4]  (.Q (read_data[4]), .CK (CTS_n_tid1_5), .D (write_data[4]));
DFF_X1 \my_reg_reg[5]  (.Q (read_data[5]), .CK (CTS_n_tid1_5), .D (write_data[5]));
DFF_X1 \my_reg_reg[6]  (.Q (read_data[6]), .CK (CTS_n_tid1_5), .D (write_data[6]));
DFF_X1 \my_reg_reg[7]  (.Q (read_data[7]), .CK (CTS_n_tid1_5), .D (write_data[7]));
DFF_X1 \my_reg_reg[8]  (.Q (read_data[8]), .CK (CTS_n_tid1_5), .D (write_data[8]));
DFF_X1 \my_reg_reg[9]  (.Q (read_data[9]), .CK (CTS_n_tid1_5), .D (write_data[9]));
DFF_X1 \my_reg_reg[10]  (.Q (read_data[10]), .CK (CTS_n_tid1_5), .D (write_data[10]));
DFF_X1 \my_reg_reg[11]  (.Q (read_data[11]), .CK (CTS_n_tid1_5), .D (write_data[11]));
DFF_X1 \my_reg_reg[12]  (.Q (read_data[12]), .CK (CTS_n_tid1_5), .D (write_data[12]));
DFF_X1 \my_reg_reg[13]  (.Q (read_data[13]), .CK (CTS_n_tid1_5), .D (write_data[13]));
DFF_X1 \my_reg_reg[14]  (.Q (read_data[14]), .CK (CTS_n_tid1_5), .D (write_data[14]));
DFF_X1 \my_reg_reg[15]  (.Q (read_data[15]), .CK (CTS_n_tid1_5), .D (write_data[15]));
DFF_X1 \my_reg_reg[16]  (.Q (read_data[16]), .CK (CTS_n_tid1_5), .D (write_data[16]));
DFF_X1 \my_reg_reg[17]  (.Q (read_data[17]), .CK (CTS_n_tid1_5), .D (write_data[17]));
DFF_X1 \my_reg_reg[18]  (.Q (read_data[18]), .CK (CTS_n_tid1_5), .D (write_data[18]));
DFF_X1 \my_reg_reg[19]  (.Q (read_data[19]), .CK (CTS_n_tid1_5), .D (write_data[19]));
DFF_X1 \my_reg_reg[20]  (.Q (read_data[20]), .CK (CTS_n_tid1_5), .D (write_data[20]));
DFF_X1 \my_reg_reg[21]  (.Q (read_data[21]), .CK (CTS_n_tid1_5), .D (write_data[21]));
DFF_X1 \my_reg_reg[22]  (.Q (read_data[22]), .CK (CTS_n_tid1_5), .D (write_data[22]));
DFF_X1 \my_reg_reg[23]  (.Q (read_data[23]), .CK (CTS_n_tid1_5), .D (write_data[23]));
DFF_X1 \my_reg_reg[24]  (.Q (read_data[24]), .CK (CTS_n_tid1_5), .D (write_data[24]));
DFF_X1 \my_reg_reg[25]  (.Q (read_data[25]), .CK (CTS_n_tid1_5), .D (write_data[25]));
DFF_X1 \my_reg_reg[26]  (.Q (read_data[26]), .CK (CTS_n_tid1_5), .D (write_data[26]));
DFF_X1 \my_reg_reg[27]  (.Q (read_data[27]), .CK (CTS_n_tid1_5), .D (write_data[27]));
DFF_X1 \my_reg_reg[28]  (.Q (read_data[28]), .CK (CTS_n_tid1_5), .D (write_data[28]));
DFF_X1 \my_reg_reg[29]  (.Q (read_data[29]), .CK (CTS_n_tid1_5), .D (write_data[29]));
DFF_X1 \my_reg_reg[30]  (.Q (read_data[30]), .CK (CTS_n_tid1_5), .D (write_data[30]));
DFF_X1 \my_reg_reg[31]  (.Q (read_data[31]), .CK (CTS_n_tid1_5), .D (write_data[31]));
DFF_X1 \my_reg2_reg[0]  (.Q (read_data2[0]), .CK (CTS_n_tid1_5), .D (write_data2[0]));
DFF_X1 \my_reg2_reg[1]  (.Q (read_data2[1]), .CK (CTS_n_tid1_5), .D (write_data2[1]));
DFF_X1 \my_reg2_reg[2]  (.Q (read_data2[2]), .CK (CTS_n_tid1_5), .D (write_data2[2]));
DFF_X1 \my_reg2_reg[3]  (.Q (read_data2[3]), .CK (CTS_n_tid1_5), .D (write_data2[3]));
DFF_X1 \my_reg2_reg[4]  (.Q (read_data2[4]), .CK (CTS_n_tid1_5), .D (write_data2[4]));
DFF_X1 \my_reg2_reg[5]  (.Q (read_data2[5]), .CK (CTS_n_tid1_5), .D (write_data2[5]));
DFF_X1 \my_reg2_reg[6]  (.Q (read_data2[6]), .CK (CTS_n_tid1_5), .D (write_data2[6]));
DFF_X1 \my_reg2_reg[7]  (.Q (read_data2[7]), .CK (CTS_n_tid1_5), .D (write_data2[7]));
DFF_X1 \my_reg2_reg[8]  (.Q (read_data2[8]), .CK (CTS_n_tid1_5), .D (write_data2[8]));
DFF_X1 \my_reg2_reg[9]  (.Q (read_data2[9]), .CK (CTS_n_tid1_5), .D (write_data2[9]));
DFF_X1 \my_reg2_reg[10]  (.Q (read_data2[10]), .CK (CTS_n_tid1_5), .D (write_data2[10]));
DFF_X1 \my_reg2_reg[11]  (.Q (read_data2[11]), .CK (CTS_n_tid1_5), .D (write_data2[11]));
DFF_X1 \my_reg2_reg[12]  (.Q (read_data2[12]), .CK (CTS_n_tid1_5), .D (write_data2[12]));
DFF_X1 \my_reg2_reg[13]  (.Q (read_data2[13]), .CK (CTS_n_tid1_5), .D (write_data2[13]));
DFF_X1 \my_reg2_reg[14]  (.Q (read_data2[14]), .CK (CTS_n_tid1_5), .D (write_data2[14]));
DFF_X1 \my_reg2_reg[15]  (.Q (read_data2[15]), .CK (CTS_n_tid1_5), .D (write_data2[15]));
DFF_X1 \my_reg2_reg[16]  (.Q (read_data2[16]), .CK (CTS_n_tid1_5), .D (write_data2[16]));
DFF_X1 \my_reg2_reg[17]  (.Q (read_data2[17]), .CK (CTS_n_tid1_5), .D (write_data2[17]));
DFF_X1 \my_reg2_reg[18]  (.Q (read_data2[18]), .CK (CTS_n_tid1_5), .D (write_data2[18]));
DFF_X1 \my_reg2_reg[19]  (.Q (read_data2[19]), .CK (CTS_n_tid1_5), .D (write_data2[19]));
DFF_X1 \my_reg2_reg[20]  (.Q (read_data2[20]), .CK (CTS_n_tid1_5), .D (write_data2[20]));
DFF_X1 \my_reg2_reg[21]  (.Q (read_data2[21]), .CK (CTS_n_tid1_5), .D (write_data2[21]));
DFF_X1 \my_reg2_reg[22]  (.Q (read_data2[22]), .CK (CTS_n_tid1_5), .D (write_data2[22]));
DFF_X1 \my_reg2_reg[23]  (.Q (read_data2[23]), .CK (CTS_n_tid1_5), .D (write_data2[23]));
DFF_X1 \my_reg2_reg[24]  (.Q (read_data2[24]), .CK (CTS_n_tid1_5), .D (write_data2[24]));
DFF_X1 \my_reg2_reg[25]  (.Q (read_data2[25]), .CK (CTS_n_tid1_5), .D (write_data2[25]));
DFF_X1 \my_reg2_reg[26]  (.Q (read_data2[26]), .CK (CTS_n_tid1_5), .D (write_data2[26]));
DFF_X1 \my_reg2_reg[27]  (.Q (read_data2[27]), .CK (CTS_n_tid1_5), .D (write_data2[27]));
DFF_X1 \my_reg2_reg[28]  (.Q (read_data2[28]), .CK (CTS_n_tid1_5), .D (write_data2[28]));
DFF_X1 \my_reg2_reg[29]  (.Q (read_data2[29]), .CK (CTS_n_tid1_5), .D (write_data2[29]));
DFF_X1 \my_reg2_reg[30]  (.Q (read_data2[30]), .CK (CTS_n_tid1_5), .D (write_data2[30]));
DFF_X1 \my_reg2_reg[31]  (.Q (read_data2[31]), .CK (CTS_n_tid1_5), .D (write_data2[31]));
CLKBUF_X3 CTS_L4_c_tid1_3 (.Z (CTS_n_tid1_5), .A (CTS_n_tid1_6));
CLKBUF_X3 CTS_L2_c_tid1_52 (.Z (clk__CTS_1_PP_0), .A (clk__CTS_1_PP_3));
CLKBUF_X1 CTS_L1_c_tid1_59 (.Z (clk__CTS_1_PP_3), .A (clk__CTS_1_PP_4));

endmodule //regFile

module Radix4 (a, b, read_data3, clk, start, start_shift, start_i);

output [63:0] read_data3;
input [31:0] a;
input [31:0] b;
input clk;
input start;
input [4:0] start_i;
input [4:0] start_shift;
wire CLOCK_slh_n313;
wire CLOCK_slh_n338;
wire CLOCK_slh_n478;
wire CLOCK_slh_n383;
wire CLOCK_slh_n473;
wire CLOCK_slh_n468;
wire CLOCK_slh_n463;
wire CLOCK_slh_n353;
wire CLOCK_slh_n458;
wire CLOCK_slh_n453;
wire CLOCK_slh_n588;
wire CLOCK_slh_n448;
wire CLOCK_slh_n438;
wire CLOCK_slh_n583;
wire CLOCK_slh_n433;
wire CLOCK_slh_n348;
wire CLOCK_slh_n308;
wire CLOCK_slh_n428;
wire CLOCK_slh_n613;
wire CLOCK_slh_n423;
wire CLOCK_slh_n343;
wire CLOCK_slh_n578;
wire CLOCK_slh_n368;
wire CLOCK_slh_n603;
wire CLOCK_slh_n418;
wire CLOCK_slh_n488;
wire CLOCK_slh_n393;
wire CLOCK_slh_n388;
wire CLOCK_slh_n483;
wire CLOCK_slh_n593;
wire CLOCK_slh_n443;
wire CLOCK_slh_n328;
wire CLOCK_slh_n363;
wire CLOCK_slh_n558;
wire CLOCK_slh_n553;
wire CLOCK_slh_n548;
wire CLOCK_slh_n358;
wire CLOCK_slh_n543;
wire CLOCK_slh_n538;
wire CLOCK_slh_n533;
wire CLOCK_slh_n528;
wire CLOCK_slh_n408;
wire CLOCK_slh_n523;
wire CLOCK_slh_n518;
wire CLOCK_slh_n513;
wire CLOCK_slh_n403;
wire CLOCK_slh_n573;
wire CLOCK_slh_n618;
wire CLOCK_slh_n508;
wire CLOCK_slh_n373;
wire CLOCK_slh_n503;
wire CLOCK_slh_n498;
wire CLOCK_slh_n398;
wire CLOCK_slh_n493;
wire CLOCK_slh_n568;
wire CLOCK_slh_n413;
wire CLOCK_slh_n563;
wire CLOCK_slh_n378;
wire CLOCK_slh_n608;
wire CLOCK_slh_n598;
wire CLOCK_slh_n333;
wire CLOCK_slh_n303;
wire CLOCK_slh_n323;
wire CLOCK_slh_n318;
wire CTS_n_tid1_147;
wire CLOCK_slh_n298;
wire \read_data2[31] ;
wire \read_data2[30] ;
wire \read_data2[29] ;
wire \read_data2[28] ;
wire \read_data2[27] ;
wire \read_data2[26] ;
wire \read_data2[25] ;
wire \read_data2[24] ;
wire \read_data2[23] ;
wire \read_data2[22] ;
wire \read_data2[21] ;
wire \read_data2[20] ;
wire \read_data2[19] ;
wire \read_data2[18] ;
wire \read_data2[17] ;
wire \read_data2[16] ;
wire \read_data2[15] ;
wire \read_data2[14] ;
wire \read_data2[13] ;
wire \read_data2[12] ;
wire \read_data2[11] ;
wire \read_data2[10] ;
wire \read_data2[9] ;
wire \read_data2[8] ;
wire \read_data2[7] ;
wire \read_data2[6] ;
wire \read_data2[5] ;
wire \read_data2[4] ;
wire \read_data2[3] ;
wire \read_data2[2] ;
wire \read_data2[1] ;
wire \read_data2[0] ;
wire \read_data[31] ;
wire \read_data[30] ;
wire \read_data[29] ;
wire \read_data[28] ;
wire \read_data[27] ;
wire \read_data[26] ;
wire \read_data[25] ;
wire \read_data[24] ;
wire \read_data[23] ;
wire \read_data[22] ;
wire \read_data[21] ;
wire \read_data[20] ;
wire \read_data[19] ;
wire \read_data[18] ;
wire \read_data[17] ;
wire \read_data[16] ;
wire \read_data[15] ;
wire \read_data[14] ;
wire \read_data[13] ;
wire \read_data[12] ;
wire \read_data[11] ;
wire \read_data[10] ;
wire \read_data[9] ;
wire \read_data[8] ;
wire \read_data[7] ;
wire \read_data[6] ;
wire \read_data[5] ;
wire \read_data[4] ;
wire \read_data[3] ;
wire \read_data[2] ;
wire \read_data[1] ;
wire \read_data[0] ;
wire CTS_n_tid0_68;
wire \res[63] ;
wire \res[62] ;
wire \res[61] ;
wire \res[60] ;
wire \res[59] ;
wire \res[58] ;
wire \res[57] ;
wire \res[56] ;
wire \res[55] ;
wire \res[54] ;
wire \res[53] ;
wire \res[52] ;
wire \res[51] ;
wire \res[50] ;
wire \res[49] ;
wire \res[48] ;
wire \res[47] ;
wire \res[46] ;
wire \res[45] ;
wire \res[44] ;
wire \res[43] ;
wire \res[42] ;
wire \res[41] ;
wire \res[40] ;
wire \res[39] ;
wire \res[38] ;
wire \res[37] ;
wire \res[36] ;
wire \res[35] ;
wire \res[34] ;
wire \res[33] ;
wire \res[32] ;
wire \res[31] ;
wire \res[30] ;
wire \res[29] ;
wire \res[28] ;
wire \res[27] ;
wire \res[26] ;
wire \res[25] ;
wire \res[24] ;
wire \res[23] ;
wire \res[22] ;
wire \res[21] ;
wire \res[20] ;
wire \res[19] ;
wire \res[18] ;
wire \res[17] ;
wire \res[16] ;
wire \res[15] ;
wire \res[14] ;
wire \res[13] ;
wire \res[12] ;
wire \res[11] ;
wire \res[10] ;
wire \res[9] ;
wire \res[8] ;
wire \res[7] ;
wire \res[6] ;
wire \res[5] ;
wire \res[4] ;
wire \res[3] ;
wire \res[2] ;
wire \res[1] ;
wire \res[0] ;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_1;
wire n_0_0_2;
wire n_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_3;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_66;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_67;
wire n_0_0_17;
wire n_0_68;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_70;
wire n_0_0_20;
wire n_0_71;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_72;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_73;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_74;
wire n_0_0_33;
wire n_0_75;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_105;
wire n_0_0_38;
wire n_0_69;
wire n_0_0_39;
wire n_0_235;
wire n_0_0_40;
wire n_0_236;
wire n_0_0_41;
wire n_0_237;
wire n_0_0_42;
wire n_0_238;
wire n_0_0_43;
wire n_0_239;
wire n_0_0_44;
wire n_0_240;
wire n_0_0_45;
wire n_0_241;
wire n_0_0_46;
wire n_0_242;
wire n_0_0_47;
wire n_0_243;
wire n_0_0_48;
wire n_0_244;
wire n_0_0_49;
wire n_0_245;
wire n_0_0_50;
wire n_0_246;
wire n_0_0_51;
wire n_0_247;
wire n_0_0_52;
wire n_0_248;
wire n_0_0_53;
wire n_0_249;
wire n_0_0_54;
wire n_0_250;
wire n_0_0_55;
wire n_0_251;
wire n_0_0_56;
wire n_0_252;
wire n_0_0_57;
wire n_0_253;
wire n_0_0_58;
wire n_0_254;
wire n_0_0_59;
wire n_0_255;
wire n_0_0_60;
wire n_0_256;
wire n_0_0_61;
wire n_0_257;
wire n_0_0_62;
wire n_0_258;
wire n_0_0_63;
wire n_0_259;
wire n_0_0_64;
wire n_0_260;
wire n_0_0_65;
wire n_0_261;
wire n_0_0_66;
wire n_0_262;
wire n_0_0_67;
wire n_0_263;
wire n_0_0_68;
wire n_0_264;
wire n_0_0_69;
wire n_0_265;
wire n_0_0_70;
wire n_0_266;
wire n_0_0_71;
wire n_0_267;
wire n_0_0_72;
wire n_0_268;
wire n_0_0_73;
wire n_0_269;
wire n_0_0_74;
wire n_0_76;
wire n_0_0_75;
wire n_0_77;
wire n_0_0_76;
wire n_0_78;
wire n_0_0_77;
wire n_0_79;
wire n_0_0_78;
wire n_0_80;
wire n_0_0_79;
wire n_0_81;
wire n_0_0_80;
wire n_0_82;
wire n_0_0_81;
wire n_0_83;
wire n_0_0_82;
wire n_0_84;
wire n_0_0_83;
wire n_0_85;
wire n_0_0_84;
wire n_0_86;
wire n_0_0_85;
wire n_0_87;
wire n_0_0_86;
wire n_0_88;
wire n_0_0_87;
wire n_0_89;
wire n_0_0_88;
wire n_0_90;
wire n_0_0_89;
wire n_0_91;
wire n_0_0_90;
wire n_0_92;
wire n_0_0_91;
wire n_0_93;
wire n_0_0_92;
wire n_0_94;
wire n_0_0_93;
wire n_0_95;
wire n_0_0_94;
wire n_0_96;
wire n_0_0_95;
wire n_0_97;
wire n_0_0_96;
wire n_0_98;
wire n_0_0_97;
wire n_0_99;
wire n_0_0_98;
wire n_0_100;
wire n_0_0_99;
wire n_0_101;
wire n_0_0_100;
wire n_0_102;
wire n_0_0_101;
wire n_0_103;
wire n_0_0_102;
wire n_0_104;
wire n_0_0_103;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_0_110;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_0_113;
wire n_0_0_114;
wire n_0_0_115;
wire n_0_0_116;
wire n_0_0_117;
wire n_0_0_118;
wire n_0_0_119;
wire n_0_0_120;
wire n_0_0_121;
wire n_0_0_122;
wire n_0_0_123;
wire n_0_0_124;
wire n_0_0_125;
wire n_0_0_126;
wire n_0_0_127;
wire n_0_0_128;
wire n_0_0_129;
wire n_0_0_130;
wire n_0_0_131;
wire n_0_0_132;
wire n_0_0_133;
wire n_0_0_134;
wire n_0_0_135;
wire n_0_0_136;
wire n_0_0_137;
wire n_0_0_138;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_144;
wire n_0_0_145;
wire n_0_0_146;
wire n_0_0_147;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_0_153;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_108;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_0_188;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_109;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_110;
wire n_0_0_207;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_111;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_112;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_0_224;
wire n_0_113;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_114;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_115;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_116;
wire n_0_0_248;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_0_253;
wire n_0_117;
wire n_0_0_254;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_118;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_119;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_0_271;
wire n_0_120;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_121;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_122;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_0_289;
wire n_0_123;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_124;
wire n_0_0_299;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_125;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_126;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_127;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_128;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_129;
wire n_0_0_339;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_130;
wire n_0_0_347;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_131;
wire n_0_0_355;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire n_0_0_360;
wire n_0_0_361;
wire n_0_0_362;
wire n_0_132;
wire n_0_0_363;
wire n_0_0_364;
wire n_0_0_365;
wire n_0_0_366;
wire n_0_0_367;
wire n_0_0_368;
wire n_0_0_369;
wire n_0_0_370;
wire n_0_0_371;
wire n_0_133;
wire n_0_0_372;
wire n_0_0_373;
wire n_0_0_374;
wire n_0_0_375;
wire n_0_0_376;
wire n_0_0_377;
wire n_0_0_378;
wire n_0_0_379;
wire n_0_134;
wire n_0_0_380;
wire n_0_0_381;
wire n_0_0_382;
wire n_0_0_383;
wire n_0_0_384;
wire n_0_0_385;
wire n_0_0_386;
wire n_0_0_387;
wire n_0_135;
wire n_0_0_388;
wire n_0_0_389;
wire n_0_0_390;
wire n_0_0_391;
wire n_0_0_392;
wire n_0_0_393;
wire n_0_0_394;
wire n_0_0_395;
wire n_0_0_396;
wire n_0_0_397;
wire n_0_136;
wire n_0_0_398;
wire n_0_0_399;
wire n_0_0_400;
wire n_0_0_401;
wire n_0_0_402;
wire n_0_0_403;
wire n_0_0_404;
wire n_0_0_405;
wire n_0_137;
wire n_0_0_406;
wire n_0_0_407;
wire n_0_0_408;
wire n_0_0_409;
wire n_0_0_410;
wire n_0_0_411;
wire n_0_0_412;
wire n_0_0_413;
wire n_0_138;
wire n_0_0_414;
wire n_0_0_415;
wire n_0_0_416;
wire n_0_0_417;
wire n_0_0_418;
wire n_0_0_419;
wire n_0_0_420;
wire n_0_0_421;
wire n_0_139;
wire n_0_0_422;
wire n_0_107;
wire n_0_0_423;
wire n_0_0_424;
wire n_0_0_425;
wire n_0_0_426;
wire n_0_0_427;
wire n_0_0_428;
wire n_0_0_429;
wire n_0_0_430;
wire n_0_0_431;
wire n_0_0_432;
wire n_0_140;
wire n_0_0_433;
wire n_0_0_434;
wire n_0_0_435;
wire n_0_0_436;
wire n_0_0_437;
wire n_0_0_438;
wire n_0_141;
wire n_0_0_439;
wire n_0_0_440;
wire n_0_0_441;
wire n_0_0_442;
wire n_0_0_443;
wire n_0_142;
wire n_0_0_444;
wire n_0_0_445;
wire n_0_0_446;
wire n_0_0_447;
wire n_0_0_448;
wire n_0_143;
wire n_0_0_449;
wire n_0_0_450;
wire n_0_0_451;
wire n_0_0_452;
wire n_0_0_453;
wire n_0_144;
wire n_0_0_454;
wire n_0_0_455;
wire n_0_0_456;
wire n_0_0_457;
wire n_0_0_458;
wire n_0_145;
wire n_0_0_459;
wire n_0_0_460;
wire n_0_0_461;
wire n_0_0_462;
wire n_0_0_463;
wire n_0_146;
wire n_0_0_464;
wire n_0_0_465;
wire n_0_0_466;
wire n_0_0_467;
wire n_0_0_468;
wire n_0_147;
wire n_0_0_469;
wire n_0_0_470;
wire n_0_0_471;
wire n_0_0_472;
wire n_0_0_473;
wire n_0_0_474;
wire n_0_148;
wire n_0_0_475;
wire n_0_0_476;
wire n_0_0_477;
wire n_0_0_478;
wire n_0_0_479;
wire n_0_0_480;
wire n_0_149;
wire n_0_0_481;
wire n_0_0_482;
wire n_0_0_483;
wire n_0_0_484;
wire n_0_0_485;
wire n_0_0_486;
wire n_0_150;
wire n_0_0_487;
wire n_0_0_488;
wire n_0_0_489;
wire n_0_0_490;
wire n_0_151;
wire n_0_0_491;
wire n_0_0_492;
wire n_0_0_493;
wire n_0_0_494;
wire n_0_0_495;
wire n_0_152;
wire n_0_0_496;
wire n_0_0_497;
wire n_0_0_498;
wire n_0_0_499;
wire n_0_153;
wire n_0_0_500;
wire n_0_0_501;
wire n_0_0_502;
wire n_0_0_503;
wire n_0_154;
wire n_0_0_504;
wire n_0_0_505;
wire n_0_0_506;
wire n_0_0_507;
wire n_0_155;
wire n_0_0_508;
wire n_0_0_509;
wire n_0_0_510;
wire n_0_0_511;
wire n_0_0_512;
wire n_0_0_513;
wire n_0_156;
wire n_0_0_514;
wire n_0_0_515;
wire n_0_0_516;
wire n_0_0_517;
wire n_0_157;
wire n_0_0_518;
wire n_0_0_519;
wire n_0_0_520;
wire n_0_0_521;
wire n_0_158;
wire n_0_0_522;
wire n_0_0_523;
wire n_0_0_524;
wire n_0_0_525;
wire n_0_159;
wire n_0_0_526;
wire n_0_0_527;
wire n_0_0_528;
wire n_0_0_529;
wire n_0_160;
wire n_0_0_530;
wire n_0_0_531;
wire n_0_0_532;
wire n_0_0_533;
wire n_0_161;
wire n_0_0_534;
wire n_0_0_535;
wire n_0_0_536;
wire n_0_0_537;
wire n_0_162;
wire n_0_0_538;
wire n_0_0_539;
wire n_0_0_540;
wire n_0_0_541;
wire n_0_163;
wire n_0_0_542;
wire n_0_0_543;
wire n_0_0_544;
wire n_0_0_545;
wire n_0_0_546;
wire n_0_164;
wire n_0_0_547;
wire n_0_0_548;
wire n_0_0_549;
wire n_0_0_550;
wire n_0_165;
wire n_0_0_551;
wire n_0_0_552;
wire n_0_0_553;
wire n_0_0_554;
wire n_0_166;
wire n_0_0_555;
wire n_0_0_556;
wire n_0_0_557;
wire n_0_0_558;
wire n_0_167;
wire n_0_0_559;
wire n_0_0_560;
wire n_0_0_561;
wire n_0_0_562;
wire n_0_0_563;
wire n_0_168;
wire n_0_0_564;
wire n_0_0_565;
wire n_0_0_566;
wire n_0_0_567;
wire n_0_169;
wire n_0_0_568;
wire n_0_0_569;
wire n_0_0_570;
wire n_0_0_571;
wire n_0_170;
wire write_en;
wire \c[63] ;
wire \c[62] ;
wire \c[61] ;
wire \c[60] ;
wire \c[59] ;
wire \c[58] ;
wire \c[57] ;
wire \c[56] ;
wire \c[55] ;
wire \c[54] ;
wire \c[53] ;
wire \c[52] ;
wire \c[51] ;
wire \c[50] ;
wire \c[49] ;
wire \c[48] ;
wire \c[47] ;
wire \c[46] ;
wire \c[45] ;
wire \c[44] ;
wire \c[43] ;
wire \c[42] ;
wire \c[41] ;
wire \c[40] ;
wire \c[39] ;
wire \c[38] ;
wire \c[37] ;
wire \c[36] ;
wire \c[35] ;
wire \c[34] ;
wire \c[33] ;
wire \c[32] ;
wire \c[31] ;
wire \c[30] ;
wire \c[29] ;
wire \c[28] ;
wire \c[27] ;
wire \c[26] ;
wire \c[25] ;
wire \c[24] ;
wire \c[23] ;
wire \c[22] ;
wire \c[21] ;
wire \c[20] ;
wire \c[19] ;
wire \c[18] ;
wire \c[17] ;
wire \c[16] ;
wire \c[15] ;
wire \c[14] ;
wire \c[13] ;
wire \c[12] ;
wire \c[11] ;
wire \c[10] ;
wire \c[9] ;
wire \c[8] ;
wire \c[7] ;
wire \c[6] ;
wire \c[5] ;
wire \c[4] ;
wire \c[3] ;
wire \c[2] ;
wire \c[1] ;
wire \c[0] ;
wire \shift[5] ;
wire \shift[4] ;
wire \shift[3] ;
wire \shift[2] ;
wire \shift[1] ;
wire \shift[0] ;
wire \i[5] ;
wire \i[4] ;
wire \i[3] ;
wire \i[2] ;
wire \i[1] ;
wire \i[0] ;
wire n_0_106;
wire uc_0;
wire uc_1;
wire uc_2;
wire hfn_ipo_n49;
wire hfn_ipo_n50;
wire hfn_ipo_n41;
wire CTS_n_tid0_69;
wire hfn_ipo_n45;
wire hfn_ipo_n46;
wire hfn_ipo_n35;
wire hfn_ipo_n36;
wire hfn_ipo_n37;
wire CTS_n_tid1_199;
wire hfn_ipo_n43;
wire hfn_ipo_n44;
wire hfn_ipo_n47;
wire hfn_ipo_n48;
wire drc_ipo_n51;
wire hfn_ipo_n39;
wire CTS_n_tid1_188;
wire CTS_n_tid1_187;
wire CLOCK_slh__n619;
wire CLOCK_slh__n621;
wire CLOCK_slh__n623;
wire CLOCK_slh__n625;
wire CLOCK_slh__n627;
wire CLOCK_slh__n629;
wire CLOCK_slh__n631;
wire CLOCK_slh__n633;
wire CLOCK_slh__n635;
wire CLOCK_slh__n637;
wire CLOCK_slh__n639;
wire CLOCK_slh__n640;
wire CLOCK_slh__n641;
wire CLOCK_slh__n645;
wire CLOCK_slh__n646;
wire CLOCK_slh__n647;
wire CLOCK_slh__n651;
wire CLOCK_slh__n652;
wire CLOCK_slh__n653;
wire CLOCK_slh__n657;
wire CLOCK_slh__n658;
wire CLOCK_slh__n659;
wire CLOCK_slh__n663;
wire CLOCK_slh__n664;
wire CLOCK_slh__n665;
wire CLOCK_slh__n669;
wire CLOCK_slh__n670;
wire CLOCK_slh__n671;
wire CLOCK_slh__n675;
wire CLOCK_slh__n676;
wire CLOCK_slh__n677;
wire CLOCK_slh__n681;
wire CLOCK_slh__n682;
wire CLOCK_slh__n683;
wire CLOCK_slh__n687;
wire CLOCK_slh__n688;
wire CLOCK_slh__n689;
wire CLOCK_slh__n693;
wire CLOCK_slh__n694;
wire CLOCK_slh__n695;
wire CLOCK_slh__n699;
wire CLOCK_slh__n700;
wire CLOCK_slh__n701;
wire CLOCK_slh__n705;
wire CLOCK_slh__n706;
wire CLOCK_slh__n707;
wire CLOCK_slh__n711;
wire CLOCK_slh__n712;
wire CLOCK_slh__n713;
wire CLOCK_slh__n717;
wire CLOCK_slh__n718;
wire CLOCK_slh__n719;
wire CLOCK_slh__n723;
wire CLOCK_slh__n724;
wire CLOCK_slh__n725;
wire CLOCK_slh__n729;
wire CLOCK_slh__n730;
wire CLOCK_slh__n731;
wire CLOCK_slh__n735;
wire CLOCK_slh__n736;
wire CLOCK_slh__n737;
wire CLOCK_slh__n741;
wire CLOCK_slh__n742;
wire CLOCK_slh__n743;
wire CLOCK_slh__n747;
wire CLOCK_slh__n748;
wire CLOCK_slh__n749;
wire CLOCK_slh__n753;
wire CLOCK_slh__n754;
wire CLOCK_slh__n755;
wire CLOCK_slh__n759;
wire CLOCK_slh__n760;
wire CLOCK_slh__n761;
wire CLOCK_slh__n765;
wire CLOCK_slh__n766;
wire CLOCK_slh__n767;
wire CLOCK_slh__n771;
wire CLOCK_slh__n772;
wire CLOCK_slh__n773;
wire CLOCK_slh__n777;
wire CLOCK_slh__n778;
wire CLOCK_slh__n779;
wire CLOCK_slh__n783;
wire CLOCK_slh__n784;
wire CLOCK_slh__n785;
wire CLOCK_slh__n789;
wire CLOCK_slh__n790;
wire CLOCK_slh__n791;
wire CLOCK_slh__n795;
wire CLOCK_slh__n796;
wire CLOCK_slh__n797;
wire CLOCK_slh__n801;
wire CLOCK_slh__n802;
wire CLOCK_slh__n803;
wire CLOCK_slh__n807;
wire CLOCK_slh__n808;
wire CLOCK_slh__n809;
wire CLOCK_slh__n813;
wire CLOCK_slh__n814;
wire CLOCK_slh__n815;
wire CLOCK_slh__n819;
wire CLOCK_slh__n820;
wire CLOCK_slh__n821;
wire CLOCK_slh__n825;
wire CLOCK_slh__n826;
wire CLOCK_slh__n827;
wire CLOCK_slh__n831;
wire CLOCK_slh__n832;
wire CLOCK_slh__n833;
wire CLOCK_slh__n837;
wire CLOCK_slh__n838;
wire CLOCK_slh__n839;
wire CLOCK_slh__n843;
wire CLOCK_slh__n844;
wire CLOCK_slh__n845;
wire CLOCK_slh__n849;
wire CLOCK_slh__n850;
wire CLOCK_slh__n851;
wire CLOCK_slh__n855;
wire CLOCK_slh__n856;
wire CLOCK_slh__n857;
wire CLOCK_slh__n861;
wire CLOCK_slh__n862;
wire CLOCK_slh__n863;
wire CLOCK_slh__n867;
wire CLOCK_slh__n868;
wire CLOCK_slh__n869;
wire CLOCK_slh__n873;
wire CLOCK_slh__n874;
wire CLOCK_slh__n875;
wire CLOCK_slh__n879;
wire CLOCK_slh__n880;
wire CLOCK_slh__n881;
wire CLOCK_slh__n885;
wire CLOCK_slh__n886;
wire CLOCK_slh__n887;
wire CLOCK_slh__n891;
wire CLOCK_slh__n892;
wire CLOCK_slh__n893;
wire CLOCK_slh__n897;
wire CLOCK_slh__n898;
wire CLOCK_slh__n899;
wire CLOCK_slh__n903;
wire CLOCK_slh__n904;
wire CLOCK_slh__n905;
wire CLOCK_slh__n909;
wire CLOCK_slh__n910;
wire CLOCK_slh__n911;
wire CLOCK_slh__n915;
wire CLOCK_slh__n916;
wire CLOCK_slh__n917;
wire CLOCK_slh__n921;
wire CLOCK_slh__n922;
wire CLOCK_slh__n923;
wire CLOCK_slh__n927;
wire CLOCK_slh__n928;
wire CLOCK_slh__n929;
wire CLOCK_slh__n933;
wire CLOCK_slh__n934;
wire CLOCK_slh__n935;
wire CLOCK_slh__n939;
wire CLOCK_slh__n940;
wire CLOCK_slh__n941;
wire CLOCK_slh__n945;
wire CLOCK_slh__n946;
wire CLOCK_slh__n947;
wire CLOCK_slh__n951;
wire CLOCK_slh__n952;
wire CLOCK_slh__n953;
wire CLOCK_slh__n957;
wire CLOCK_slh__n958;
wire CLOCK_slh__n959;
wire CLOCK_slh__n963;
wire CLOCK_slh__n964;
wire CLOCK_slh__n965;
wire CLOCK_slh__n969;
wire CLOCK_slh__n970;
wire CLOCK_slh__n971;
wire CLOCK_slh__n975;
wire CLOCK_slh__n976;
wire CLOCK_slh__n977;
wire CLOCK_slh__n981;
wire CLOCK_slh__n982;
wire CLOCK_slh__n983;
wire CLOCK_slh__n987;
wire CLOCK_slh__n988;
wire CLOCK_slh__n989;
wire CLOCK_slh__n993;
wire CLOCK_slh__n994;
wire CLOCK_slh__n995;
wire CLOCK_slh__n999;
wire CLOCK_slh__n1000;
wire CLOCK_slh__n1001;
wire CLOCK_slh__n1005;
wire CLOCK_slh__n1006;
wire CLOCK_slh__n1007;
wire CLOCK_slh__n1011;
wire CLOCK_slh__n1012;
wire CLOCK_slh__n1013;
wire CLOCK_slh__n1017;
wire CLOCK_slh__n1018;
wire CLOCK_slh__n1019;


CLKGATETST_X1 clk_gate_i_reg (.GCK (n_0_106), .CK (CTS_n_tid1_188), .E (n_0_69), .SE (1'b0 ));
DFF_X1 \i_reg[0]  (.Q (\i[0] ), .CK (n_0_106), .D (n_0_1));
DFF_X1 \i_reg[1]  (.Q (\i[1] ), .CK (n_0_106), .D (n_0_2));
DFF_X1 \i_reg[2]  (.Q (\i[2] ), .CK (n_0_106), .D (n_0_3));
DFF_X1 \i_reg[3]  (.Q (\i[3] ), .CK (n_0_106), .D (n_0_66));
DFF_X1 \i_reg[4]  (.Q (\i[4] ), .CK (n_0_106), .D (n_0_67));
DFF_X1 \i_reg[5]  (.Q (\i[5] ), .CK (n_0_106), .D (n_0_68));
DFF_X1 \shift_reg[0]  (.Q (\shift[0] ), .CK (n_0_106), .D (n_0_70));
DFF_X1 \shift_reg[1]  (.Q (\shift[1] ), .CK (n_0_106), .D (n_0_71));
DFF_X1 \shift_reg[2]  (.Q (\shift[2] ), .CK (n_0_106), .D (n_0_72));
DFF_X1 \shift_reg[3]  (.Q (\shift[3] ), .CK (n_0_106), .D (n_0_73));
DFF_X1 \shift_reg[4]  (.Q (\shift[4] ), .CK (n_0_106), .D (n_0_74));
DFF_X1 \shift_reg[5]  (.Q (\shift[5] ), .CK (n_0_106), .D (n_0_75));
DFF_X1 \c_reg[0]  (.Q (\c[0] ), .CK (CTS_n_tid1_147), .D (n_0_235));
DFF_X1 \c_reg[1]  (.Q (\c[1] ), .CK (CTS_n_tid1_147), .D (n_0_236));
DFF_X1 \c_reg[2]  (.Q (\c[2] ), .CK (CTS_n_tid1_147), .D (n_0_237));
DFF_X1 \c_reg[3]  (.Q (\c[3] ), .CK (CTS_n_tid1_147), .D (n_0_238));
DFF_X1 \c_reg[4]  (.Q (\c[4] ), .CK (CTS_n_tid1_147), .D (n_0_239));
DFF_X1 \c_reg[5]  (.Q (\c[5] ), .CK (CTS_n_tid1_147), .D (n_0_240));
DFF_X1 \c_reg[6]  (.Q (\c[6] ), .CK (CTS_n_tid1_147), .D (n_0_241));
DFF_X1 \c_reg[7]  (.Q (\c[7] ), .CK (CTS_n_tid1_147), .D (n_0_242));
DFF_X1 \c_reg[8]  (.Q (\c[8] ), .CK (CTS_n_tid1_147), .D (n_0_243));
DFF_X1 \c_reg[9]  (.Q (\c[9] ), .CK (CTS_n_tid1_147), .D (n_0_244));
DFF_X1 \c_reg[10]  (.Q (\c[10] ), .CK (CTS_n_tid1_147), .D (n_0_245));
DFF_X1 \c_reg[11]  (.Q (\c[11] ), .CK (CTS_n_tid1_147), .D (n_0_246));
DFF_X1 \c_reg[12]  (.Q (\c[12] ), .CK (CTS_n_tid1_147), .D (n_0_247));
DFF_X1 \c_reg[13]  (.Q (\c[13] ), .CK (CTS_n_tid1_147), .D (n_0_248));
DFF_X1 \c_reg[14]  (.Q (\c[14] ), .CK (CTS_n_tid1_147), .D (n_0_249));
DFF_X1 \c_reg[15]  (.Q (\c[15] ), .CK (CTS_n_tid1_147), .D (n_0_250));
DFF_X1 \c_reg[16]  (.Q (\c[16] ), .CK (CTS_n_tid1_147), .D (n_0_251));
DFF_X1 \c_reg[17]  (.Q (\c[17] ), .CK (CTS_n_tid1_147), .D (n_0_252));
DFF_X1 \c_reg[18]  (.Q (\c[18] ), .CK (CTS_n_tid1_147), .D (n_0_253));
DFF_X1 \c_reg[19]  (.Q (\c[19] ), .CK (CTS_n_tid1_147), .D (n_0_254));
DFF_X1 \c_reg[20]  (.Q (\c[20] ), .CK (CTS_n_tid1_147), .D (n_0_255));
DFF_X1 \c_reg[21]  (.Q (\c[21] ), .CK (CTS_n_tid1_147), .D (n_0_256));
DFF_X1 \c_reg[22]  (.Q (\c[22] ), .CK (CTS_n_tid1_147), .D (n_0_257));
DFF_X1 \c_reg[23]  (.Q (\c[23] ), .CK (CTS_n_tid1_147), .D (n_0_258));
DFF_X1 \c_reg[24]  (.Q (\c[24] ), .CK (CTS_n_tid1_147), .D (n_0_259));
DFF_X1 \c_reg[25]  (.Q (\c[25] ), .CK (CTS_n_tid1_147), .D (n_0_260));
DFF_X1 \c_reg[26]  (.Q (\c[26] ), .CK (CTS_n_tid1_187), .D (n_0_261));
DFF_X1 \c_reg[27]  (.Q (\c[27] ), .CK (CTS_n_tid1_187), .D (n_0_262));
DFF_X1 \c_reg[28]  (.Q (\c[28] ), .CK (CTS_n_tid1_187), .D (n_0_263));
DFF_X1 \c_reg[29]  (.Q (\c[29] ), .CK (CTS_n_tid1_187), .D (n_0_264));
DFF_X1 \c_reg[30]  (.Q (\c[30] ), .CK (CTS_n_tid1_187), .D (n_0_265));
DFF_X1 \c_reg[31]  (.Q (\c[31] ), .CK (CTS_n_tid1_187), .D (n_0_266));
DFF_X1 \c_reg[32]  (.Q (\c[32] ), .CK (CTS_n_tid1_187), .D (n_0_267));
DFF_X1 \c_reg[33]  (.Q (\c[33] ), .CK (CTS_n_tid1_187), .D (n_0_268));
DFF_X1 \c_reg[34]  (.Q (\c[34] ), .CK (CTS_n_tid1_187), .D (n_0_269));
DFF_X1 \c_reg[35]  (.Q (\c[35] ), .CK (CTS_n_tid1_187), .D (n_0_76));
DFF_X1 \c_reg[36]  (.Q (\c[36] ), .CK (CTS_n_tid1_187), .D (n_0_77));
DFF_X1 \c_reg[37]  (.Q (\c[37] ), .CK (CTS_n_tid1_187), .D (n_0_78));
DFF_X1 \c_reg[38]  (.Q (\c[38] ), .CK (CTS_n_tid1_187), .D (n_0_79));
DFF_X1 \c_reg[39]  (.Q (\c[39] ), .CK (CTS_n_tid1_187), .D (n_0_80));
DFF_X1 \c_reg[40]  (.Q (\c[40] ), .CK (CTS_n_tid1_187), .D (n_0_81));
DFF_X1 \c_reg[41]  (.Q (\c[41] ), .CK (CTS_n_tid1_187), .D (n_0_82));
DFF_X1 \c_reg[42]  (.Q (\c[42] ), .CK (CTS_n_tid1_187), .D (n_0_83));
DFF_X1 \c_reg[43]  (.Q (\c[43] ), .CK (CTS_n_tid1_187), .D (n_0_84));
DFF_X1 \c_reg[44]  (.Q (\c[44] ), .CK (CTS_n_tid1_187), .D (n_0_85));
DFF_X1 \c_reg[45]  (.Q (\c[45] ), .CK (CTS_n_tid1_187), .D (n_0_86));
DFF_X1 \c_reg[46]  (.Q (\c[46] ), .CK (CTS_n_tid1_187), .D (n_0_87));
DFF_X1 \c_reg[47]  (.Q (\c[47] ), .CK (CTS_n_tid1_187), .D (n_0_88));
DFF_X1 \c_reg[48]  (.Q (\c[48] ), .CK (CTS_n_tid1_187), .D (n_0_89));
DFF_X1 \c_reg[49]  (.Q (\c[49] ), .CK (CTS_n_tid1_187), .D (n_0_90));
DFF_X1 \c_reg[50]  (.Q (\c[50] ), .CK (CTS_n_tid1_187), .D (n_0_91));
DFF_X1 \c_reg[51]  (.Q (\c[51] ), .CK (CTS_n_tid1_187), .D (n_0_92));
DFF_X1 \c_reg[52]  (.Q (\c[52] ), .CK (CTS_n_tid1_187), .D (n_0_93));
DFF_X1 \c_reg[53]  (.Q (\c[53] ), .CK (CTS_n_tid1_187), .D (n_0_94));
DFF_X1 \c_reg[54]  (.Q (\c[54] ), .CK (CTS_n_tid1_187), .D (n_0_95));
DFF_X1 \c_reg[55]  (.Q (\c[55] ), .CK (CTS_n_tid1_187), .D (n_0_96));
DFF_X1 \c_reg[56]  (.Q (\c[56] ), .CK (CTS_n_tid1_187), .D (n_0_97));
DFF_X1 \c_reg[57]  (.Q (\c[57] ), .CK (CTS_n_tid1_187), .D (n_0_98));
DFF_X1 \c_reg[58]  (.Q (\c[58] ), .CK (CTS_n_tid1_187), .D (n_0_99));
DFF_X1 \c_reg[59]  (.Q (\c[59] ), .CK (CTS_n_tid1_187), .D (n_0_100));
DFF_X1 \c_reg[60]  (.Q (\c[60] ), .CK (CTS_n_tid1_187), .D (n_0_101));
DFF_X1 \c_reg[61]  (.Q (\c[61] ), .CK (CTS_n_tid1_187), .D (n_0_102));
DFF_X1 \c_reg[62]  (.Q (\c[62] ), .CK (CTS_n_tid1_187), .D (n_0_103));
DFF_X1 \c_reg[63]  (.Q (\c[63] ), .CK (CTS_n_tid1_187), .D (n_0_104));
DFF_X1 write_en_reg (.Q (write_en), .CK (CTS_n_tid1_147), .D (CLOCK_slh_n298));
OAI21_X1 i_0_0_713 (.ZN (n_0_170), .A (n_0_0_571), .B1 (hfn_ipo_n36), .B2 (n_0_0_567));
OAI221_X1 i_0_0_712 (.ZN (n_0_0_571), .A (hfn_ipo_n36), .B1 (hfn_ipo_n48), .B2 (n_0_0_570)
    , .C1 (n_0_0_562), .C2 (n_0_0_24));
OAI22_X1 i_0_0_711 (.ZN (n_0_0_570), .A1 (n_0_0_552), .A2 (n_0_0_23), .B1 (n_0_0_568), .B2 (n_0_0_569));
AOI21_X1 i_0_0_710 (.ZN (n_0_0_569), .A (n_0_0_509), .B1 (n_0_0_410), .B2 (\shift[5] ));
OAI21_X1 i_0_0_709 (.ZN (n_0_0_568), .A (n_0_0_23), .B1 (n_0_0_534), .B2 (n_0_0_543));
OAI22_X1 i_0_0_708 (.ZN (n_0_169), .A1 (n_0_0_563), .A2 (hfn_ipo_n36), .B1 (n_0_0_567), .B2 (hfn_ipo_n50));
OAI22_X1 i_0_0_707 (.ZN (n_0_0_567), .A1 (n_0_0_557), .A2 (n_0_0_24), .B1 (hfn_ipo_n48), .B2 (n_0_0_566));
OAI22_X1 i_0_0_706 (.ZN (n_0_0_566), .A1 (n_0_0_548), .A2 (n_0_0_23), .B1 (n_0_0_564), .B2 (n_0_0_565));
AOI21_X1 i_0_0_705 (.ZN (n_0_0_565), .A (n_0_0_509), .B1 (n_0_0_402), .B2 (\shift[5] ));
OAI21_X1 i_0_0_704 (.ZN (n_0_0_564), .A (n_0_0_23), .B1 (n_0_0_530), .B2 (n_0_0_543));
OAI22_X1 i_0_0_703 (.ZN (n_0_168), .A1 (n_0_0_563), .A2 (hfn_ipo_n50), .B1 (n_0_0_558), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_702 (.ZN (n_0_0_563), .A1 (n_0_0_562), .A2 (n_0_0_24), .B1 (n_0_0_553), .B2 (hfn_ipo_n48));
OAI21_X1 i_0_0_701 (.ZN (n_0_0_562), .A (n_0_0_561), .B1 (n_0_0_23), .B2 (n_0_0_544));
OAI211_X1 i_0_0_700 (.ZN (n_0_0_561), .A (n_0_0_560), .B (hfn_ipo_n37), .C1 (n_0_0_526), .C2 (n_0_0_543));
OAI221_X1 i_0_0_699 (.ZN (n_0_0_560), .A (n_0_0_295), .B1 (n_0_0_392), .B2 (n_0_0_428)
    , .C1 (n_0_0_491), .C2 (n_0_0_559));
INV_X1 i_0_0_698 (.ZN (n_0_0_559), .A (n_0_0_428));
OAI22_X1 i_0_0_697 (.ZN (n_0_167), .A1 (n_0_0_558), .A2 (hfn_ipo_n50), .B1 (n_0_0_554), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_696 (.ZN (n_0_0_558), .A1 (n_0_0_557), .A2 (n_0_0_24), .B1 (n_0_0_549), .B2 (hfn_ipo_n48));
AOI22_X1 i_0_0_695 (.ZN (n_0_0_557), .A1 (n_0_0_539), .A2 (hfn_ipo_n46), .B1 (n_0_0_556), .B2 (n_0_0_23));
AOI221_X1 i_0_0_694 (.ZN (n_0_0_556), .A (n_0_0_423), .B1 (n_0_0_384), .B2 (n_0_0_555)
    , .C1 (\shift[3] ), .C2 (n_0_0_522));
NOR2_X1 i_0_0_693 (.ZN (n_0_0_555), .A1 (n_0_0_33), .A2 (\shift[3] ));
OAI22_X1 i_0_0_692 (.ZN (n_0_166), .A1 (n_0_0_550), .A2 (hfn_ipo_n36), .B1 (n_0_0_554), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_691 (.ZN (n_0_0_554), .A1 (n_0_0_553), .A2 (n_0_0_24), .B1 (n_0_0_545), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_690 (.ZN (n_0_0_553), .A1 (n_0_0_535), .A2 (n_0_0_23), .B1 (hfn_ipo_n46), .B2 (n_0_0_552));
OAI22_X1 i_0_0_689 (.ZN (n_0_0_552), .A1 (n_0_0_551), .A2 (n_0_0_509), .B1 (n_0_0_518), .B2 (n_0_0_543));
NOR2_X1 i_0_0_688 (.ZN (n_0_0_551), .A1 (n_0_0_375), .A2 (n_0_0_33));
OAI22_X1 i_0_0_687 (.ZN (n_0_165), .A1 (n_0_0_546), .A2 (hfn_ipo_n36), .B1 (n_0_0_550), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_686 (.ZN (n_0_0_550), .A1 (n_0_0_540), .A2 (hfn_ipo_n48), .B1 (n_0_0_549), .B2 (n_0_0_24));
OAI22_X1 i_0_0_685 (.ZN (n_0_0_549), .A1 (n_0_0_531), .A2 (n_0_0_23), .B1 (hfn_ipo_n46), .B2 (n_0_0_548));
OAI22_X1 i_0_0_684 (.ZN (n_0_0_548), .A1 (n_0_0_547), .A2 (n_0_0_509), .B1 (n_0_0_514), .B2 (n_0_0_543));
NOR2_X1 i_0_0_683 (.ZN (n_0_0_547), .A1 (n_0_0_367), .A2 (n_0_0_33));
OAI22_X1 i_0_0_682 (.ZN (n_0_164), .A1 (n_0_0_541), .A2 (hfn_ipo_n36), .B1 (n_0_0_546), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_681 (.ZN (n_0_0_546), .A1 (n_0_0_536), .A2 (hfn_ipo_n48), .B1 (n_0_0_24), .B2 (n_0_0_545));
OAI22_X1 i_0_0_680 (.ZN (n_0_0_545), .A1 (n_0_0_527), .A2 (n_0_0_23), .B1 (hfn_ipo_n46), .B2 (n_0_0_544));
OAI22_X1 i_0_0_679 (.ZN (n_0_0_544), .A1 (n_0_0_542), .A2 (n_0_0_509), .B1 (n_0_0_510), .B2 (n_0_0_543));
NAND2_X1 i_0_0_678 (.ZN (n_0_0_543), .A1 (n_0_0_424), .A2 (\shift[3] ));
NOR2_X1 i_0_0_677 (.ZN (n_0_0_542), .A1 (n_0_0_358), .A2 (n_0_0_33));
OAI22_X1 i_0_0_676 (.ZN (n_0_163), .A1 (n_0_0_541), .A2 (hfn_ipo_n50), .B1 (n_0_0_537), .B2 (hfn_ipo_n36));
OAI22_X1 i_0_0_675 (.ZN (n_0_0_541), .A1 (n_0_0_532), .A2 (n_0_0_24), .B1 (n_0_0_540), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_674 (.ZN (n_0_0_540), .A1 (n_0_0_523), .A2 (n_0_0_23), .B1 (n_0_0_539), .B2 (hfn_ipo_n46));
OAI21_X1 i_0_0_673 (.ZN (n_0_0_539), .A (n_0_0_538), .B1 (n_0_0_504), .B2 (n_0_0_295));
OAI21_X1 i_0_0_672 (.ZN (n_0_0_538), .A (n_0_0_508), .B1 (n_0_0_33), .B2 (n_0_0_350));
OAI22_X1 i_0_0_671 (.ZN (n_0_162), .A1 (n_0_0_533), .A2 (hfn_ipo_n36), .B1 (n_0_0_537), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_670 (.ZN (n_0_0_537), .A1 (n_0_0_536), .A2 (n_0_0_24), .B1 (n_0_0_528), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_669 (.ZN (n_0_0_536), .A1 (n_0_0_519), .A2 (n_0_0_23), .B1 (n_0_0_535), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_668 (.ZN (n_0_0_535), .A1 (n_0_0_500), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_534));
NOR2_X1 i_0_0_667 (.ZN (n_0_0_534), .A1 (n_0_0_342), .A2 (n_0_0_33));
OAI22_X1 i_0_0_666 (.ZN (n_0_161), .A1 (n_0_0_533), .A2 (hfn_ipo_n50), .B1 (n_0_0_529), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_665 (.ZN (n_0_0_533), .A1 (n_0_0_524), .A2 (hfn_ipo_n48), .B1 (n_0_0_532), .B2 (n_0_0_24));
AOI22_X1 i_0_0_664 (.ZN (n_0_0_532), .A1 (n_0_0_515), .A2 (hfn_ipo_n46), .B1 (n_0_0_531), .B2 (n_0_0_23));
OAI22_X1 i_0_0_663 (.ZN (n_0_0_531), .A1 (n_0_0_496), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_530));
NOR2_X1 i_0_0_662 (.ZN (n_0_0_530), .A1 (n_0_0_334), .A2 (n_0_0_33));
OAI22_X1 i_0_0_661 (.ZN (n_0_160), .A1 (n_0_0_525), .A2 (hfn_ipo_n36), .B1 (n_0_0_529), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_660 (.ZN (n_0_0_529), .A1 (n_0_0_520), .A2 (hfn_ipo_n48), .B1 (n_0_0_528), .B2 (n_0_0_24));
OAI22_X1 i_0_0_659 (.ZN (n_0_0_528), .A1 (n_0_0_511), .A2 (n_0_0_23), .B1 (n_0_0_527), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_658 (.ZN (n_0_0_527), .A1 (n_0_0_492), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_526));
NOR2_X1 i_0_0_657 (.ZN (n_0_0_526), .A1 (n_0_0_326), .A2 (n_0_0_33));
OAI22_X1 i_0_0_656 (.ZN (n_0_159), .A1 (n_0_0_525), .A2 (hfn_ipo_n50), .B1 (n_0_0_521), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_655 (.ZN (n_0_0_525), .A1 (n_0_0_516), .A2 (hfn_ipo_n48), .B1 (n_0_0_524), .B2 (n_0_0_24));
OAI22_X1 i_0_0_654 (.ZN (n_0_0_524), .A1 (n_0_0_505), .A2 (n_0_0_23), .B1 (n_0_0_523), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_653 (.ZN (n_0_0_523), .A1 (n_0_0_487), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_522));
NOR2_X1 i_0_0_652 (.ZN (n_0_0_522), .A1 (n_0_0_318), .A2 (n_0_0_33));
OAI22_X1 i_0_0_651 (.ZN (n_0_158), .A1 (n_0_0_517), .A2 (hfn_ipo_n36), .B1 (n_0_0_521), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_650 (.ZN (n_0_0_521), .A1 (n_0_0_520), .A2 (n_0_0_24), .B1 (n_0_0_512), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_649 (.ZN (n_0_0_520), .A1 (n_0_0_501), .A2 (n_0_0_23), .B1 (n_0_0_519), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_648 (.ZN (n_0_0_519), .A1 (n_0_0_483), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_518));
NOR2_X1 i_0_0_647 (.ZN (n_0_0_518), .A1 (n_0_0_310), .A2 (n_0_0_33));
OAI22_X1 i_0_0_646 (.ZN (n_0_157), .A1 (n_0_0_517), .A2 (hfn_ipo_n50), .B1 (n_0_0_513), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_645 (.ZN (n_0_0_517), .A1 (hfn_ipo_n48), .A2 (n_0_0_506), .B1 (n_0_0_516), .B2 (n_0_0_24));
OAI22_X1 i_0_0_644 (.ZN (n_0_0_516), .A1 (n_0_0_497), .A2 (n_0_0_23), .B1 (n_0_0_515), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_643 (.ZN (n_0_0_515), .A1 (n_0_0_477), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_514));
NOR2_X1 i_0_0_642 (.ZN (n_0_0_514), .A1 (n_0_0_302), .A2 (n_0_0_33));
OAI22_X1 i_0_0_641 (.ZN (n_0_156), .A1 (n_0_0_507), .A2 (hfn_ipo_n36), .B1 (n_0_0_513), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_640 (.ZN (n_0_0_513), .A1 (n_0_0_502), .A2 (hfn_ipo_n48), .B1 (n_0_0_512), .B2 (n_0_0_24));
OAI22_X1 i_0_0_639 (.ZN (n_0_0_512), .A1 (n_0_0_511), .A2 (hfn_ipo_n46), .B1 (n_0_0_493), .B2 (n_0_0_23));
OAI22_X1 i_0_0_638 (.ZN (n_0_0_511), .A1 (n_0_0_471), .A2 (n_0_0_295), .B1 (n_0_0_509), .B2 (n_0_0_510));
NOR2_X1 i_0_0_637 (.ZN (n_0_0_510), .A1 (n_0_0_293), .A2 (n_0_0_33));
INV_X1 i_0_0_636 (.ZN (n_0_0_509), .A (n_0_0_508));
NOR2_X1 i_0_0_635 (.ZN (n_0_0_508), .A1 (n_0_0_423), .A2 (\shift[3] ));
OAI22_X1 i_0_0_634 (.ZN (n_0_155), .A1 (n_0_0_507), .A2 (hfn_ipo_n50), .B1 (n_0_0_503), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_633 (.ZN (n_0_0_507), .A1 (n_0_0_498), .A2 (hfn_ipo_n48), .B1 (n_0_0_506), .B2 (n_0_0_24));
OAI22_X1 i_0_0_632 (.ZN (n_0_0_506), .A1 (n_0_0_505), .A2 (hfn_ipo_n46), .B1 (n_0_0_488), .B2 (n_0_0_23));
AOI22_X1 i_0_0_631 (.ZN (n_0_0_505), .A1 (n_0_0_465), .A2 (\shift[3] ), .B1 (n_0_0_504), .B2 (n_0_0_295));
OAI221_X1 i_0_0_630 (.ZN (n_0_0_504), .A (n_0_0_433), .B1 (n_0_0_417), .B2 (n_0_0_428)
    , .C1 (n_0_0_389), .C2 (n_0_0_416));
OAI22_X1 i_0_0_629 (.ZN (n_0_154), .A1 (n_0_0_499), .A2 (hfn_ipo_n36), .B1 (n_0_0_503), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_628 (.ZN (n_0_0_503), .A1 (n_0_0_502), .A2 (n_0_0_24), .B1 (n_0_0_494), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_627 (.ZN (n_0_0_502), .A1 (n_0_0_484), .A2 (n_0_0_23), .B1 (n_0_0_501), .B2 (hfn_ipo_n46));
AOI22_X1 i_0_0_626 (.ZN (n_0_0_501), .A1 (n_0_0_460), .A2 (\shift[3] ), .B1 (n_0_0_500), .B2 (n_0_0_295));
OAI221_X1 i_0_0_625 (.ZN (n_0_0_500), .A (n_0_0_433), .B1 (n_0_0_406), .B2 (n_0_0_428)
    , .C1 (n_0_0_389), .C2 (n_0_0_409));
OAI22_X1 i_0_0_624 (.ZN (n_0_153), .A1 (n_0_0_499), .A2 (hfn_ipo_n50), .B1 (n_0_0_495), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_623 (.ZN (n_0_0_499), .A1 (n_0_0_498), .A2 (n_0_0_24), .B1 (n_0_0_489), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_622 (.ZN (n_0_0_498), .A1 (n_0_0_497), .A2 (hfn_ipo_n46), .B1 (n_0_0_478), .B2 (n_0_0_23));
AOI22_X1 i_0_0_621 (.ZN (n_0_0_497), .A1 (n_0_0_455), .A2 (\shift[3] ), .B1 (n_0_0_496), .B2 (n_0_0_295));
OAI221_X1 i_0_0_620 (.ZN (n_0_0_496), .A (n_0_0_433), .B1 (n_0_0_398), .B2 (n_0_0_428)
    , .C1 (n_0_0_389), .C2 (n_0_0_401));
OAI22_X1 i_0_0_619 (.ZN (n_0_152), .A1 (n_0_0_490), .A2 (hfn_ipo_n36), .B1 (n_0_0_495), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_618 (.ZN (n_0_0_495), .A1 (n_0_0_485), .A2 (hfn_ipo_n48), .B1 (n_0_0_494), .B2 (n_0_0_24));
OAI22_X1 i_0_0_617 (.ZN (n_0_0_494), .A1 (n_0_0_493), .A2 (hfn_ipo_n46), .B1 (n_0_0_472), .B2 (n_0_0_23));
AOI22_X1 i_0_0_616 (.ZN (n_0_0_493), .A1 (n_0_0_450), .A2 (\shift[3] ), .B1 (n_0_0_492), .B2 (n_0_0_295));
OAI22_X1 i_0_0_615 (.ZN (n_0_0_492), .A1 (n_0_0_491), .A2 (\shift[4] ), .B1 (n_0_0_389), .B2 (n_0_0_392));
AOI21_X1 i_0_0_614 (.ZN (n_0_0_491), .A (n_0_0_423), .B1 (\shift[5] ), .B2 (n_0_0_268));
OAI22_X1 i_0_0_613 (.ZN (n_0_151), .A1 (n_0_0_490), .A2 (hfn_ipo_n50), .B1 (n_0_0_486), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_612 (.ZN (n_0_0_490), .A1 (n_0_0_479), .A2 (hfn_ipo_n48), .B1 (n_0_0_489), .B2 (n_0_0_24));
OAI22_X1 i_0_0_611 (.ZN (n_0_0_489), .A1 (n_0_0_488), .A2 (hfn_ipo_n46), .B1 (n_0_0_466), .B2 (n_0_0_23));
OAI22_X1 i_0_0_610 (.ZN (n_0_0_488), .A1 (n_0_0_445), .A2 (n_0_0_295), .B1 (n_0_0_487), .B2 (\shift[3] ));
OAI221_X1 i_0_0_609 (.ZN (n_0_0_487), .A (n_0_0_433), .B1 (n_0_0_383), .B2 (n_0_0_389)
    , .C1 (n_0_0_380), .C2 (n_0_0_428));
OAI22_X1 i_0_0_608 (.ZN (n_0_150), .A1 (n_0_0_480), .A2 (hfn_ipo_n36), .B1 (n_0_0_486), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_607 (.ZN (n_0_0_486), .A1 (n_0_0_485), .A2 (n_0_0_24), .B1 (n_0_0_473), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_606 (.ZN (n_0_0_485), .A1 (n_0_0_484), .A2 (hfn_ipo_n46), .B1 (n_0_0_461), .B2 (n_0_0_23));
AOI22_X1 i_0_0_605 (.ZN (n_0_0_484), .A1 (n_0_0_440), .A2 (\shift[3] ), .B1 (n_0_0_483), .B2 (n_0_0_295));
OAI221_X1 i_0_0_604 (.ZN (n_0_0_483), .A (n_0_0_433), .B1 (n_0_0_481), .B2 (n_0_0_428)
    , .C1 (n_0_0_482), .C2 (n_0_0_389));
INV_X1 i_0_0_603 (.ZN (n_0_0_482), .A (n_0_0_374));
INV_X1 i_0_0_602 (.ZN (n_0_0_481), .A (n_0_0_256));
OAI22_X1 i_0_0_601 (.ZN (n_0_149), .A1 (n_0_0_480), .A2 (hfn_ipo_n50), .B1 (n_0_0_474), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_600 (.ZN (n_0_0_480), .A1 (n_0_0_479), .A2 (n_0_0_24), .B1 (n_0_0_467), .B2 (hfn_ipo_n48));
AOI22_X1 i_0_0_599 (.ZN (n_0_0_479), .A1 (n_0_0_478), .A2 (n_0_0_23), .B1 (n_0_0_456), .B2 (hfn_ipo_n46));
OAI22_X1 i_0_0_598 (.ZN (n_0_0_478), .A1 (n_0_0_477), .A2 (\shift[3] ), .B1 (n_0_0_435), .B2 (n_0_0_295));
OAI221_X1 i_0_0_597 (.ZN (n_0_0_477), .A (n_0_0_433), .B1 (n_0_0_475), .B2 (n_0_0_389)
    , .C1 (n_0_0_476), .C2 (n_0_0_428));
INV_X1 i_0_0_596 (.ZN (n_0_0_476), .A (n_0_0_250));
INV_X1 i_0_0_595 (.ZN (n_0_0_475), .A (n_0_0_366));
OAI22_X1 i_0_0_594 (.ZN (n_0_148), .A1 (n_0_0_468), .A2 (hfn_ipo_n36), .B1 (n_0_0_474), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_593 (.ZN (n_0_0_474), .A1 (n_0_0_462), .A2 (hfn_ipo_n48), .B1 (n_0_0_473), .B2 (n_0_0_24));
OAI22_X1 i_0_0_592 (.ZN (n_0_0_473), .A1 (n_0_0_451), .A2 (n_0_0_23), .B1 (n_0_0_472), .B2 (hfn_ipo_n46));
AOI22_X1 i_0_0_591 (.ZN (n_0_0_472), .A1 (n_0_0_471), .A2 (n_0_0_295), .B1 (n_0_0_429), .B2 (\shift[3] ));
OAI221_X1 i_0_0_590 (.ZN (n_0_0_471), .A (n_0_0_433), .B1 (n_0_0_469), .B2 (n_0_0_428)
    , .C1 (n_0_0_470), .C2 (n_0_0_389));
INV_X1 i_0_0_589 (.ZN (n_0_0_470), .A (n_0_0_357));
INV_X1 i_0_0_588 (.ZN (n_0_0_469), .A (n_0_0_241));
OAI22_X1 i_0_0_587 (.ZN (n_0_147), .A1 (n_0_0_468), .A2 (hfn_ipo_n50), .B1 (n_0_0_463), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_586 (.ZN (n_0_0_468), .A1 (n_0_0_457), .A2 (hfn_ipo_n48), .B1 (n_0_0_467), .B2 (n_0_0_24));
OAI22_X1 i_0_0_585 (.ZN (n_0_0_467), .A1 (n_0_0_466), .A2 (hfn_ipo_n46), .B1 (n_0_0_446), .B2 (n_0_0_23));
AOI22_X1 i_0_0_584 (.ZN (n_0_0_466), .A1 (n_0_0_465), .A2 (n_0_0_295), .B1 (\shift[3] ), .B2 (n_0_0_418));
OAI221_X1 i_0_0_583 (.ZN (n_0_0_465), .A (n_0_0_433), .B1 (n_0_0_464), .B2 (n_0_0_389)
    , .C1 (n_0_0_235), .C2 (n_0_0_428));
INV_X1 i_0_0_582 (.ZN (n_0_0_464), .A (n_0_0_349));
OAI22_X1 i_0_0_581 (.ZN (n_0_146), .A1 (n_0_0_463), .A2 (hfn_ipo_n50), .B1 (n_0_0_458), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_580 (.ZN (n_0_0_463), .A1 (n_0_0_462), .A2 (n_0_0_24), .B1 (n_0_0_452), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_579 (.ZN (n_0_0_462), .A1 (n_0_0_461), .A2 (hfn_ipo_n46), .B1 (n_0_0_441), .B2 (n_0_0_23));
AOI22_X1 i_0_0_578 (.ZN (n_0_0_461), .A1 (n_0_0_460), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_410));
OAI221_X1 i_0_0_577 (.ZN (n_0_0_460), .A (n_0_0_433), .B1 (n_0_0_229), .B2 (n_0_0_428)
    , .C1 (n_0_0_459), .C2 (n_0_0_389));
INV_X1 i_0_0_576 (.ZN (n_0_0_459), .A (n_0_0_341));
OAI22_X1 i_0_0_575 (.ZN (n_0_145), .A1 (n_0_0_458), .A2 (hfn_ipo_n50), .B1 (n_0_0_453), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_574 (.ZN (n_0_0_458), .A1 (n_0_0_457), .A2 (n_0_0_24), .B1 (n_0_0_447), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_573 (.ZN (n_0_0_457), .A1 (n_0_0_436), .A2 (n_0_0_23), .B1 (n_0_0_456), .B2 (hfn_ipo_n46));
AOI22_X1 i_0_0_572 (.ZN (n_0_0_456), .A1 (n_0_0_455), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_402));
OAI221_X1 i_0_0_571 (.ZN (n_0_0_455), .A (n_0_0_433), .B1 (n_0_0_222), .B2 (n_0_0_428)
    , .C1 (n_0_0_454), .C2 (n_0_0_389));
INV_X1 i_0_0_570 (.ZN (n_0_0_454), .A (n_0_0_333));
OAI22_X1 i_0_0_569 (.ZN (n_0_144), .A1 (n_0_0_448), .A2 (hfn_ipo_n36), .B1 (n_0_0_453), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_568 (.ZN (n_0_0_453), .A1 (n_0_0_452), .A2 (n_0_0_24), .B1 (n_0_0_442), .B2 (hfn_ipo_n48));
OAI22_X1 i_0_0_567 (.ZN (n_0_0_452), .A1 (n_0_0_451), .A2 (hfn_ipo_n46), .B1 (hfn_ipo_n37), .B2 (n_0_0_430));
AOI22_X1 i_0_0_566 (.ZN (n_0_0_451), .A1 (n_0_0_450), .A2 (n_0_0_295), .B1 (\shift[3] ), .B2 (n_0_0_394));
OAI221_X1 i_0_0_565 (.ZN (n_0_0_450), .A (n_0_0_433), .B1 (n_0_0_215), .B2 (n_0_0_428)
    , .C1 (n_0_0_449), .C2 (n_0_0_389));
INV_X1 i_0_0_564 (.ZN (n_0_0_449), .A (n_0_0_325));
OAI22_X1 i_0_0_563 (.ZN (n_0_143), .A1 (n_0_0_448), .A2 (hfn_ipo_n50), .B1 (n_0_0_443), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_562 (.ZN (n_0_0_448), .A1 (n_0_0_437), .A2 (hfn_ipo_n48), .B1 (n_0_0_447), .B2 (n_0_0_24));
OAI22_X1 i_0_0_561 (.ZN (n_0_0_447), .A1 (n_0_0_446), .A2 (hfn_ipo_n46), .B1 (hfn_ipo_n37), .B2 (n_0_0_419));
AOI22_X1 i_0_0_560 (.ZN (n_0_0_446), .A1 (n_0_0_445), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_384));
OAI221_X1 i_0_0_559 (.ZN (n_0_0_445), .A (n_0_0_433), .B1 (n_0_0_236), .B2 (n_0_0_428)
    , .C1 (n_0_0_444), .C2 (n_0_0_389));
INV_X1 i_0_0_558 (.ZN (n_0_0_444), .A (n_0_0_317));
OAI22_X1 i_0_0_557 (.ZN (n_0_142), .A1 (n_0_0_443), .A2 (hfn_ipo_n50), .B1 (n_0_0_438), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_0_556 (.ZN (n_0_0_443), .A1 (n_0_0_442), .A2 (n_0_0_24), .B1 (hfn_ipo_n48), .B2 (n_0_0_431));
OAI22_X1 i_0_0_555 (.ZN (n_0_0_442), .A1 (n_0_0_441), .A2 (hfn_ipo_n46), .B1 (hfn_ipo_n37), .B2 (n_0_0_411));
AOI22_X1 i_0_0_554 (.ZN (n_0_0_441), .A1 (n_0_0_440), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_376));
OAI221_X1 i_0_0_553 (.ZN (n_0_0_440), .A (n_0_0_433), .B1 (n_0_0_225), .B2 (n_0_0_428)
    , .C1 (n_0_0_439), .C2 (n_0_0_389));
INV_X1 i_0_0_552 (.ZN (n_0_0_439), .A (n_0_0_309));
OAI22_X1 i_0_0_551 (.ZN (n_0_141), .A1 (n_0_0_438), .A2 (hfn_ipo_n50), .B1 (hfn_ipo_n36), .B2 (n_0_0_432));
AOI22_X1 i_0_0_550 (.ZN (n_0_0_438), .A1 (n_0_0_437), .A2 (n_0_0_24), .B1 (hfn_ipo_n48), .B2 (n_0_0_420));
OAI22_X1 i_0_0_549 (.ZN (n_0_0_437), .A1 (n_0_0_436), .A2 (hfn_ipo_n46), .B1 (hfn_ipo_n37), .B2 (n_0_0_403));
AOI22_X1 i_0_0_548 (.ZN (n_0_0_436), .A1 (n_0_0_435), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_368));
OAI221_X1 i_0_0_547 (.ZN (n_0_0_435), .A (n_0_0_433), .B1 (n_0_0_434), .B2 (n_0_0_389)
    , .C1 (n_0_0_198), .C2 (n_0_0_428));
INV_X1 i_0_0_546 (.ZN (n_0_0_434), .A (n_0_0_301));
INV_X1 i_0_0_545 (.ZN (n_0_0_433), .A (n_0_0_425));
OAI22_X1 i_0_0_544 (.ZN (n_0_140), .A1 (n_0_0_432), .A2 (hfn_ipo_n50), .B1 (n_0_0_421), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_543 (.ZN (n_0_0_432), .A1 (n_0_0_431), .A2 (hfn_ipo_n39), .B1 (hfn_ipo_n47), .B2 (n_0_0_412));
OAI22_X1 i_0_0_542 (.ZN (n_0_0_431), .A1 (n_0_0_430), .A2 (hfn_ipo_n45), .B1 (hfn_ipo_n37), .B2 (n_0_0_395));
AOI22_X1 i_0_0_541 (.ZN (n_0_0_430), .A1 (n_0_0_429), .A2 (n_0_0_295), .B1 (n_0_0_363), .B2 (n_0_0_359));
OAI21_X1 i_0_0_540 (.ZN (n_0_0_429), .A (n_0_0_427), .B1 (n_0_0_171), .B2 (n_0_0_428));
NAND2_X1 i_0_0_539 (.ZN (n_0_0_428), .A1 (n_0_0_173), .A2 (\shift[5] ));
AOI21_X1 i_0_0_538 (.ZN (n_0_0_427), .A (n_0_0_425), .B1 (n_0_0_292), .B2 (n_0_0_426));
INV_X1 i_0_0_537 (.ZN (n_0_0_426), .A (n_0_0_389));
NOR2_X1 i_0_0_536 (.ZN (n_0_0_425), .A1 (n_0_0_424), .A2 (\shift[4] ));
INV_X1 i_0_0_535 (.ZN (n_0_0_424), .A (n_0_0_423));
AND2_X1 i_0_0_534 (.ZN (n_0_0_423), .A1 (n_0_107), .A2 (n_0_0_33));
NAND2_X1 i_0_0_533 (.ZN (n_0_107), .A1 (n_0_0_414), .A2 (n_0_0_422));
AOI22_X1 i_0_0_532 (.ZN (n_0_0_422), .A1 (n_0_0_200), .A2 (n_0_65), .B1 (\read_data2[31] ), .B2 (drc_ipo_n51));
OAI22_X1 i_0_0_531 (.ZN (n_0_139), .A1 (n_0_0_421), .A2 (hfn_ipo_n50), .B1 (n_0_0_413), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_530 (.ZN (n_0_0_421), .A1 (n_0_0_404), .A2 (hfn_ipo_n47), .B1 (n_0_0_420), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_529 (.ZN (n_0_0_420), .A1 (n_0_0_385), .A2 (hfn_ipo_n37), .B1 (n_0_0_419), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_528 (.ZN (n_0_0_419), .A1 (n_0_0_418), .A2 (n_0_0_295), .B1 (n_0_0_351), .B2 (n_0_0_363));
OAI22_X1 i_0_0_527 (.ZN (n_0_0_418), .A1 (n_0_0_416), .A2 (n_0_0_393), .B1 (n_0_0_417), .B2 (n_0_0_389));
INV_X1 i_0_0_526 (.ZN (n_0_0_417), .A (n_0_0_286));
AND2_X1 i_0_0_525 (.ZN (n_0_0_416), .A1 (n_0_0_414), .A2 (n_0_0_415));
AOI22_X1 i_0_0_524 (.ZN (n_0_0_415), .A1 (n_0_0_200), .A2 (n_0_64), .B1 (\read_data2[30] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_523 (.ZN (n_0_0_414), .A1 (n_0_0_196), .A2 (n_0_34), .B1 (n_0_0_197), .B2 (\read_data2[31] ));
OAI22_X1 i_0_0_522 (.ZN (n_0_138), .A1 (n_0_0_405), .A2 (hfn_ipo_n35), .B1 (n_0_0_413), .B2 (hfn_ipo_n50));
AOI22_X1 i_0_0_521 (.ZN (n_0_0_413), .A1 (n_0_0_396), .A2 (hfn_ipo_n47), .B1 (n_0_0_412), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_520 (.ZN (n_0_0_412), .A1 (n_0_0_377), .A2 (hfn_ipo_n37), .B1 (n_0_0_411), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_519 (.ZN (n_0_0_411), .A1 (n_0_0_343), .A2 (n_0_0_363), .B1 (n_0_0_410), .B2 (n_0_0_172));
OAI22_X1 i_0_0_518 (.ZN (n_0_0_410), .A1 (n_0_0_406), .A2 (n_0_0_173), .B1 (n_0_0_409), .B2 (\shift[4] ));
AND2_X1 i_0_0_517 (.ZN (n_0_0_409), .A1 (n_0_0_407), .A2 (n_0_0_408));
AOI22_X1 i_0_0_516 (.ZN (n_0_0_408), .A1 (n_0_0_197), .A2 (\read_data2[30] ), .B1 (\read_data2[29] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_515 (.ZN (n_0_0_407), .A1 (n_0_0_196), .A2 (n_0_33), .B1 (n_0_0_200), .B2 (n_0_63));
INV_X1 i_0_0_514 (.ZN (n_0_0_406), .A (n_0_0_280));
OAI22_X1 i_0_0_513 (.ZN (n_0_137), .A1 (n_0_0_405), .A2 (hfn_ipo_n49), .B1 (n_0_0_397), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_512 (.ZN (n_0_0_405), .A1 (n_0_0_404), .A2 (hfn_ipo_n39), .B1 (n_0_0_386), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_511 (.ZN (n_0_0_404), .A1 (n_0_0_369), .A2 (hfn_ipo_n37), .B1 (n_0_0_403), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_510 (.ZN (n_0_0_403), .A1 (n_0_0_335), .A2 (n_0_0_363), .B1 (n_0_0_402), .B2 (n_0_0_172));
OAI22_X1 i_0_0_509 (.ZN (n_0_0_402), .A1 (n_0_0_398), .A2 (n_0_0_173), .B1 (n_0_0_401), .B2 (\shift[4] ));
AND2_X1 i_0_0_508 (.ZN (n_0_0_401), .A1 (n_0_0_399), .A2 (n_0_0_400));
AOI22_X1 i_0_0_507 (.ZN (n_0_0_400), .A1 (n_0_0_196), .A2 (n_0_32), .B1 (\read_data2[28] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_506 (.ZN (n_0_0_399), .A1 (n_0_0_197), .A2 (\read_data2[29] ), .B1 (n_0_0_200), .B2 (n_0_62));
INV_X1 i_0_0_505 (.ZN (n_0_0_398), .A (n_0_0_274));
OAI22_X1 i_0_0_504 (.ZN (n_0_136), .A1 (n_0_0_387), .A2 (hfn_ipo_n35), .B1 (n_0_0_397), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_503 (.ZN (n_0_0_397), .A1 (n_0_0_396), .A2 (hfn_ipo_n39), .B1 (n_0_0_378), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_502 (.ZN (n_0_0_396), .A1 (n_0_0_395), .A2 (hfn_ipo_n45), .B1 (n_0_0_360), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_501 (.ZN (n_0_0_395), .A1 (n_0_0_394), .A2 (n_0_0_295), .B1 (n_0_0_327), .B2 (n_0_0_363));
OAI22_X1 i_0_0_500 (.ZN (n_0_0_394), .A1 (n_0_0_388), .A2 (n_0_0_389), .B1 (n_0_0_392), .B2 (n_0_0_393));
NAND2_X1 i_0_0_499 (.ZN (n_0_0_393), .A1 (n_0_0_173), .A2 (n_0_0_33));
AND2_X1 i_0_0_498 (.ZN (n_0_0_392), .A1 (n_0_0_390), .A2 (n_0_0_391));
AOI22_X1 i_0_0_497 (.ZN (n_0_0_391), .A1 (n_0_0_196), .A2 (n_0_31), .B1 (\read_data2[27] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_496 (.ZN (n_0_0_390), .A1 (n_0_0_197), .A2 (\read_data2[28] ), .B1 (n_0_0_200), .B2 (n_0_61));
NAND2_X1 i_0_0_495 (.ZN (n_0_0_389), .A1 (n_0_0_33), .A2 (\shift[4] ));
INV_X1 i_0_0_494 (.ZN (n_0_0_388), .A (n_0_0_268));
OAI22_X1 i_0_0_493 (.ZN (n_0_135), .A1 (n_0_0_387), .A2 (hfn_ipo_n49), .B1 (n_0_0_379), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_492 (.ZN (n_0_0_387), .A1 (n_0_0_370), .A2 (hfn_ipo_n47), .B1 (n_0_0_386), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_491 (.ZN (n_0_0_386), .A1 (n_0_0_385), .A2 (hfn_ipo_n45), .B1 (n_0_0_352), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_490 (.ZN (n_0_0_385), .A1 (n_0_0_319), .A2 (\shift[3] ), .B1 (n_0_0_384), .B2 (n_0_0_172));
AOI22_X1 i_0_0_489 (.ZN (n_0_0_384), .A1 (n_0_0_380), .A2 (\shift[4] ), .B1 (n_0_0_383), .B2 (n_0_0_173));
AND2_X1 i_0_0_488 (.ZN (n_0_0_383), .A1 (n_0_0_381), .A2 (n_0_0_382));
AOI22_X1 i_0_0_487 (.ZN (n_0_0_382), .A1 (n_0_0_197), .A2 (\read_data2[27] ), .B1 (\read_data2[26] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_486 (.ZN (n_0_0_381), .A1 (n_0_0_196), .A2 (n_0_30), .B1 (n_0_0_200), .B2 (n_0_60));
INV_X1 i_0_0_485 (.ZN (n_0_0_380), .A (n_0_0_262));
OAI22_X1 i_0_0_484 (.ZN (n_0_134), .A1 (n_0_0_379), .A2 (hfn_ipo_n49), .B1 (n_0_0_371), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_483 (.ZN (n_0_0_379), .A1 (n_0_0_361), .A2 (hfn_ipo_n47), .B1 (n_0_0_378), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_482 (.ZN (n_0_0_378), .A1 (n_0_0_377), .A2 (hfn_ipo_n45), .B1 (n_0_0_344), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_481 (.ZN (n_0_0_377), .A1 (n_0_0_311), .A2 (n_0_0_363), .B1 (n_0_0_376), .B2 (n_0_0_172));
INV_X1 i_0_0_480 (.ZN (n_0_0_376), .A (n_0_0_375));
OAI22_X1 i_0_0_479 (.ZN (n_0_0_375), .A1 (n_0_0_374), .A2 (\shift[4] ), .B1 (n_0_0_256), .B2 (n_0_0_173));
NAND2_X1 i_0_0_478 (.ZN (n_0_0_374), .A1 (n_0_0_372), .A2 (n_0_0_373));
AOI22_X1 i_0_0_477 (.ZN (n_0_0_373), .A1 (n_0_0_197), .A2 (\read_data2[26] ), .B1 (\read_data2[25] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_476 (.ZN (n_0_0_372), .A1 (n_0_0_196), .A2 (n_0_29), .B1 (n_0_0_200), .B2 (n_0_59));
OAI22_X1 i_0_0_475 (.ZN (n_0_133), .A1 (n_0_0_362), .A2 (hfn_ipo_n35), .B1 (n_0_0_371), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_474 (.ZN (n_0_0_371), .A1 (n_0_0_370), .A2 (hfn_ipo_n39), .B1 (n_0_0_353), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_473 (.ZN (n_0_0_370), .A1 (n_0_0_369), .A2 (hfn_ipo_n45), .B1 (n_0_0_336), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_472 (.ZN (n_0_0_369), .A1 (n_0_0_303), .A2 (n_0_0_363), .B1 (n_0_0_368), .B2 (n_0_0_172));
INV_X1 i_0_0_471 (.ZN (n_0_0_368), .A (n_0_0_367));
OAI22_X1 i_0_0_470 (.ZN (n_0_0_367), .A1 (n_0_0_250), .A2 (n_0_0_173), .B1 (n_0_0_366), .B2 (\shift[4] ));
NAND2_X1 i_0_0_469 (.ZN (n_0_0_366), .A1 (n_0_0_364), .A2 (n_0_0_365));
AOI22_X1 i_0_0_468 (.ZN (n_0_0_365), .A1 (n_0_0_196), .A2 (n_0_28), .B1 (\read_data2[24] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_467 (.ZN (n_0_0_364), .A1 (n_0_0_197), .A2 (\read_data2[25] ), .B1 (n_0_0_200), .B2 (n_0_58));
INV_X1 i_0_0_466 (.ZN (n_0_0_363), .A (n_0_0_243));
OAI22_X1 i_0_0_465 (.ZN (n_0_132), .A1 (n_0_0_362), .A2 (hfn_ipo_n49), .B1 (n_0_0_354), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_464 (.ZN (n_0_0_362), .A1 (n_0_0_361), .A2 (hfn_ipo_n39), .B1 (n_0_0_345), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_463 (.ZN (n_0_0_361), .A1 (n_0_0_360), .A2 (hfn_ipo_n45), .B1 (n_0_0_328), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_462 (.ZN (n_0_0_360), .A1 (n_0_0_294), .A2 (\shift[3] ), .B1 (n_0_0_359), .B2 (n_0_0_172));
INV_X1 i_0_0_461 (.ZN (n_0_0_359), .A (n_0_0_358));
AOI22_X1 i_0_0_460 (.ZN (n_0_0_358), .A1 (n_0_0_357), .A2 (n_0_0_173), .B1 (n_0_0_241), .B2 (\shift[4] ));
NAND2_X1 i_0_0_459 (.ZN (n_0_0_357), .A1 (n_0_0_355), .A2 (n_0_0_356));
AOI22_X1 i_0_0_458 (.ZN (n_0_0_356), .A1 (n_0_0_197), .A2 (\read_data2[24] ), .B1 (\read_data2[23] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_457 (.ZN (n_0_0_355), .A1 (n_0_0_196), .A2 (n_0_27), .B1 (n_0_0_200), .B2 (n_0_57));
OAI22_X1 i_0_0_456 (.ZN (n_0_131), .A1 (n_0_0_346), .A2 (hfn_ipo_n35), .B1 (n_0_0_354), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_455 (.ZN (n_0_0_354), .A1 (n_0_0_337), .A2 (hfn_ipo_n47), .B1 (n_0_0_353), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_454 (.ZN (n_0_0_353), .A1 (n_0_0_352), .A2 (hfn_ipo_n45), .B1 (n_0_0_320), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_453 (.ZN (n_0_0_352), .A1 (n_0_0_351), .A2 (n_0_0_172), .B1 (n_0_0_286), .B2 (n_0_0_244));
INV_X1 i_0_0_452 (.ZN (n_0_0_351), .A (n_0_0_350));
OAI22_X1 i_0_0_451 (.ZN (n_0_0_350), .A1 (n_0_0_349), .A2 (\shift[4] ), .B1 (n_0_0_234), .B2 (n_0_0_173));
NAND2_X1 i_0_0_450 (.ZN (n_0_0_349), .A1 (n_0_0_347), .A2 (n_0_0_348));
AOI22_X1 i_0_0_449 (.ZN (n_0_0_348), .A1 (n_0_0_196), .A2 (n_0_26), .B1 (\read_data2[22] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_448 (.ZN (n_0_0_347), .A1 (n_0_0_197), .A2 (\read_data2[23] ), .B1 (n_0_0_200), .B2 (n_0_56));
OAI22_X1 i_0_0_447 (.ZN (n_0_130), .A1 (n_0_0_346), .A2 (hfn_ipo_n49), .B1 (n_0_0_338), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_446 (.ZN (n_0_0_346), .A1 (n_0_0_329), .A2 (hfn_ipo_n47), .B1 (n_0_0_345), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_445 (.ZN (n_0_0_345), .A1 (n_0_0_312), .A2 (hfn_ipo_n37), .B1 (n_0_0_344), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_444 (.ZN (n_0_0_344), .A1 (n_0_0_343), .A2 (n_0_0_172), .B1 (n_0_0_280), .B2 (n_0_0_244));
INV_X1 i_0_0_443 (.ZN (n_0_0_343), .A (n_0_0_342));
OAI22_X1 i_0_0_442 (.ZN (n_0_0_342), .A1 (n_0_0_228), .A2 (n_0_0_173), .B1 (n_0_0_341), .B2 (\shift[4] ));
NAND2_X1 i_0_0_441 (.ZN (n_0_0_341), .A1 (n_0_0_339), .A2 (n_0_0_340));
AOI22_X1 i_0_0_440 (.ZN (n_0_0_340), .A1 (n_0_0_196), .A2 (n_0_25), .B1 (\read_data2[21] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_439 (.ZN (n_0_0_339), .A1 (n_0_0_197), .A2 (\read_data2[22] ), .B1 (n_0_0_200), .B2 (n_0_55));
OAI22_X1 i_0_0_438 (.ZN (n_0_129), .A1 (n_0_0_338), .A2 (hfn_ipo_n49), .B1 (n_0_0_330), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_437 (.ZN (n_0_0_338), .A1 (n_0_0_337), .A2 (hfn_ipo_n39), .B1 (n_0_0_321), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_436 (.ZN (n_0_0_337), .A1 (n_0_0_304), .A2 (hfn_ipo_n37), .B1 (n_0_0_336), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_435 (.ZN (n_0_0_336), .A1 (n_0_0_335), .A2 (n_0_0_172), .B1 (n_0_0_274), .B2 (n_0_0_244));
INV_X1 i_0_0_434 (.ZN (n_0_0_335), .A (n_0_0_334));
OAI22_X1 i_0_0_433 (.ZN (n_0_0_334), .A1 (n_0_0_221), .A2 (n_0_0_173), .B1 (n_0_0_333), .B2 (\shift[4] ));
NAND2_X1 i_0_0_432 (.ZN (n_0_0_333), .A1 (n_0_0_331), .A2 (n_0_0_332));
AOI22_X1 i_0_0_431 (.ZN (n_0_0_332), .A1 (n_0_0_196), .A2 (n_0_24), .B1 (\read_data2[20] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_430 (.ZN (n_0_0_331), .A1 (n_0_0_197), .A2 (\read_data2[21] ), .B1 (n_0_0_200), .B2 (n_0_54));
OAI22_X1 i_0_0_429 (.ZN (n_0_128), .A1 (hfn_ipo_n49), .A2 (n_0_0_330), .B1 (n_0_0_322), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_428 (.ZN (n_0_0_330), .A1 (n_0_0_329), .A2 (hfn_ipo_n39), .B1 (n_0_0_313), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_427 (.ZN (n_0_0_329), .A1 (n_0_0_328), .A2 (hfn_ipo_n45), .B1 (n_0_0_296), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_426 (.ZN (n_0_0_328), .A1 (n_0_0_327), .A2 (n_0_0_172), .B1 (n_0_0_268), .B2 (n_0_0_244));
INV_X1 i_0_0_425 (.ZN (n_0_0_327), .A (n_0_0_326));
OAI22_X1 i_0_0_424 (.ZN (n_0_0_326), .A1 (n_0_0_214), .A2 (n_0_0_173), .B1 (n_0_0_325), .B2 (\shift[4] ));
NAND2_X1 i_0_0_423 (.ZN (n_0_0_325), .A1 (n_0_0_323), .A2 (n_0_0_324));
AOI22_X1 i_0_0_422 (.ZN (n_0_0_324), .A1 (n_0_0_196), .A2 (n_0_23), .B1 (\read_data2[19] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_421 (.ZN (n_0_0_323), .A1 (n_0_0_197), .A2 (\read_data2[20] ), .B1 (n_0_0_200), .B2 (n_0_53));
OAI22_X1 i_0_0_420 (.ZN (n_0_127), .A1 (hfn_ipo_n35), .A2 (n_0_0_314), .B1 (n_0_0_322), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_419 (.ZN (n_0_0_322), .A1 (n_0_0_305), .A2 (hfn_ipo_n47), .B1 (n_0_0_321), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_418 (.ZN (n_0_0_321), .A1 (n_0_0_320), .A2 (hfn_ipo_n45), .B1 (hfn_ipo_n37), .B2 (n_0_0_287));
AOI22_X1 i_0_0_417 (.ZN (n_0_0_320), .A1 (n_0_0_319), .A2 (n_0_0_295), .B1 (n_0_0_262), .B2 (n_0_0_244));
NOR2_X1 i_0_0_416 (.ZN (n_0_0_319), .A1 (n_0_0_318), .A2 (\shift[5] ));
OAI22_X1 i_0_0_415 (.ZN (n_0_0_318), .A1 (n_0_0_209), .A2 (n_0_0_173), .B1 (n_0_0_317), .B2 (\shift[4] ));
NAND2_X1 i_0_0_414 (.ZN (n_0_0_317), .A1 (n_0_0_315), .A2 (n_0_0_316));
AOI22_X1 i_0_0_413 (.ZN (n_0_0_316), .A1 (n_0_0_196), .A2 (n_0_22), .B1 (\read_data2[18] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_412 (.ZN (n_0_0_315), .A1 (n_0_0_197), .A2 (\read_data2[19] ), .B1 (n_0_0_200), .B2 (n_0_52));
OAI22_X1 i_0_0_411 (.ZN (n_0_126), .A1 (n_0_0_314), .A2 (hfn_ipo_n49), .B1 (n_0_0_306), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_410 (.ZN (n_0_0_314), .A1 (n_0_0_297), .A2 (hfn_ipo_n47), .B1 (n_0_0_313), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_409 (.ZN (n_0_0_313), .A1 (n_0_0_312), .A2 (hfn_ipo_n45), .B1 (hfn_ipo_n37), .B2 (n_0_0_281));
AOI22_X1 i_0_0_408 (.ZN (n_0_0_312), .A1 (n_0_0_311), .A2 (n_0_0_172), .B1 (n_0_0_256), .B2 (n_0_0_244));
INV_X1 i_0_0_407 (.ZN (n_0_0_311), .A (n_0_0_310));
OAI22_X1 i_0_0_406 (.ZN (n_0_0_310), .A1 (n_0_0_203), .A2 (n_0_0_173), .B1 (n_0_0_309), .B2 (\shift[4] ));
NAND2_X1 i_0_0_405 (.ZN (n_0_0_309), .A1 (n_0_0_307), .A2 (n_0_0_308));
AOI22_X1 i_0_0_404 (.ZN (n_0_0_308), .A1 (n_0_0_196), .A2 (n_0_21), .B1 (\read_data2[17] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_403 (.ZN (n_0_0_307), .A1 (n_0_0_197), .A2 (\read_data2[18] ), .B1 (n_0_0_200), .B2 (n_0_51));
OAI22_X1 i_0_0_402 (.ZN (n_0_125), .A1 (n_0_0_306), .A2 (hfn_ipo_n49), .B1 (n_0_0_298), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_401 (.ZN (n_0_0_306), .A1 (n_0_0_305), .A2 (hfn_ipo_n39), .B1 (hfn_ipo_n47), .B2 (n_0_0_288));
OAI22_X1 i_0_0_400 (.ZN (n_0_0_305), .A1 (n_0_0_304), .A2 (hfn_ipo_n45), .B1 (hfn_ipo_n37), .B2 (n_0_0_275));
AOI22_X1 i_0_0_399 (.ZN (n_0_0_304), .A1 (n_0_0_303), .A2 (n_0_0_172), .B1 (n_0_0_244), .B2 (n_0_0_250));
INV_X1 i_0_0_398 (.ZN (n_0_0_303), .A (n_0_0_302));
OAI22_X1 i_0_0_397 (.ZN (n_0_0_302), .A1 (n_0_0_301), .A2 (\shift[4] ), .B1 (n_0_0_210), .B2 (n_0_0_173));
NAND2_X1 i_0_0_396 (.ZN (n_0_0_301), .A1 (n_0_0_299), .A2 (n_0_0_300));
AOI22_X1 i_0_0_395 (.ZN (n_0_0_300), .A1 (n_0_0_197), .A2 (\read_data2[17] ), .B1 (\read_data2[16] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_394 (.ZN (n_0_0_299), .A1 (n_0_0_196), .A2 (n_0_20), .B1 (n_0_0_200), .B2 (n_0_50));
OAI22_X1 i_0_0_393 (.ZN (n_0_124), .A1 (n_0_0_298), .A2 (hfn_ipo_n49), .B1 (hfn_ipo_n35), .B2 (n_0_0_289));
AOI22_X1 i_0_0_392 (.ZN (n_0_0_298), .A1 (n_0_0_297), .A2 (hfn_ipo_n39), .B1 (hfn_ipo_n47), .B2 (n_0_0_282));
OAI22_X1 i_0_0_391 (.ZN (n_0_0_297), .A1 (n_0_0_296), .A2 (hfn_ipo_n45), .B1 (hfn_ipo_n37), .B2 (n_0_0_269));
AOI22_X1 i_0_0_390 (.ZN (n_0_0_296), .A1 (n_0_0_294), .A2 (n_0_0_295), .B1 (n_0_0_241), .B2 (n_0_0_244));
INV_X1 i_0_0_389 (.ZN (n_0_0_295), .A (\shift[3] ));
NOR2_X1 i_0_0_388 (.ZN (n_0_0_294), .A1 (n_0_0_293), .A2 (\shift[5] ));
AOI22_X1 i_0_0_387 (.ZN (n_0_0_293), .A1 (n_0_0_292), .A2 (n_0_0_173), .B1 (\shift[4] ), .B2 (n_0_0_204));
NAND2_X1 i_0_0_386 (.ZN (n_0_0_292), .A1 (n_0_0_290), .A2 (n_0_0_291));
AOI22_X1 i_0_0_385 (.ZN (n_0_0_291), .A1 (n_0_0_197), .A2 (\read_data2[16] ), .B1 (\read_data2[15] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_384 (.ZN (n_0_0_290), .A1 (n_0_0_196), .A2 (n_0_19), .B1 (n_0_0_200), .B2 (n_0_49));
OAI22_X1 i_0_0_383 (.ZN (n_0_123), .A1 (n_0_0_289), .A2 (hfn_ipo_n49), .B1 (n_0_0_283), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_382 (.ZN (n_0_0_289), .A1 (n_0_0_288), .A2 (hfn_ipo_n39), .B1 (n_0_0_276), .B2 (hfn_ipo_n47));
AOI22_X1 i_0_0_381 (.ZN (n_0_0_288), .A1 (n_0_0_263), .A2 (hfn_ipo_n45), .B1 (n_0_0_287), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_380 (.ZN (n_0_0_287), .A1 (n_0_0_234), .A2 (n_0_0_244), .B1 (n_0_0_286), .B2 (n_0_0_242));
NAND2_X1 i_0_0_379 (.ZN (n_0_0_286), .A1 (n_0_0_284), .A2 (n_0_0_285));
AOI22_X1 i_0_0_378 (.ZN (n_0_0_285), .A1 (n_0_0_197), .A2 (\read_data2[15] ), .B1 (\read_data2[14] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_377 (.ZN (n_0_0_284), .A1 (n_0_0_196), .A2 (n_0_18), .B1 (n_0_0_200), .B2 (n_0_48));
OAI22_X1 i_0_0_376 (.ZN (n_0_122), .A1 (n_0_0_277), .A2 (hfn_ipo_n35), .B1 (n_0_0_283), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_375 (.ZN (n_0_0_283), .A1 (n_0_0_282), .A2 (hfn_ipo_n39), .B1 (n_0_0_270), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_374 (.ZN (n_0_0_282), .A1 (n_0_0_257), .A2 (hfn_ipo_n37), .B1 (n_0_0_281), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_373 (.ZN (n_0_0_281), .A1 (n_0_0_280), .A2 (n_0_0_242), .B1 (n_0_0_228), .B2 (n_0_0_244));
NAND2_X1 i_0_0_372 (.ZN (n_0_0_280), .A1 (n_0_0_278), .A2 (n_0_0_279));
AOI22_X1 i_0_0_371 (.ZN (n_0_0_279), .A1 (n_0_0_197), .A2 (\read_data2[14] ), .B1 (\read_data2[13] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_370 (.ZN (n_0_0_278), .A1 (n_0_0_196), .A2 (n_0_17), .B1 (n_0_0_200), .B2 (n_0_47));
OAI22_X1 i_0_0_369 (.ZN (n_0_121), .A1 (n_0_0_277), .A2 (hfn_ipo_n49), .B1 (n_0_0_271), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_368 (.ZN (n_0_0_277), .A1 (n_0_0_276), .A2 (hfn_ipo_n39), .B1 (n_0_0_264), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_367 (.ZN (n_0_0_276), .A1 (n_0_0_251), .A2 (hfn_ipo_n37), .B1 (n_0_0_275), .B2 (hfn_ipo_n45));
AOI22_X1 i_0_0_366 (.ZN (n_0_0_275), .A1 (n_0_0_221), .A2 (n_0_0_244), .B1 (n_0_0_274), .B2 (n_0_0_242));
NAND2_X1 i_0_0_365 (.ZN (n_0_0_274), .A1 (n_0_0_272), .A2 (n_0_0_273));
AOI22_X1 i_0_0_364 (.ZN (n_0_0_273), .A1 (n_0_0_196), .A2 (n_0_16), .B1 (\read_data2[12] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_363 (.ZN (n_0_0_272), .A1 (n_0_0_197), .A2 (\read_data2[13] ), .B1 (n_0_0_200), .B2 (n_0_46));
OAI22_X1 i_0_0_362 (.ZN (n_0_120), .A1 (n_0_0_265), .A2 (hfn_ipo_n35), .B1 (n_0_0_271), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_361 (.ZN (n_0_0_271), .A1 (n_0_0_270), .A2 (hfn_ipo_n39), .B1 (n_0_0_258), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_360 (.ZN (n_0_0_270), .A1 (n_0_0_269), .A2 (hfn_ipo_n45), .B1 (n_0_0_245), .B2 (hfn_ipo_n37));
AOI22_X1 i_0_0_359 (.ZN (n_0_0_269), .A1 (n_0_0_268), .A2 (n_0_0_242), .B1 (n_0_0_214), .B2 (n_0_0_244));
NAND2_X1 i_0_0_358 (.ZN (n_0_0_268), .A1 (n_0_0_266), .A2 (n_0_0_267));
AOI22_X1 i_0_0_357 (.ZN (n_0_0_267), .A1 (n_0_0_200), .A2 (n_0_45), .B1 (\read_data2[11] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_356 (.ZN (n_0_0_266), .A1 (n_0_0_197), .A2 (\read_data2[12] ), .B1 (n_0_0_196), .B2 (n_0_15));
OAI22_X1 i_0_0_355 (.ZN (n_0_119), .A1 (n_0_0_265), .A2 (hfn_ipo_n49), .B1 (n_0_0_259), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_354 (.ZN (n_0_0_265), .A1 (n_0_0_264), .A2 (hfn_ipo_n39), .B1 (n_0_0_252), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_353 (.ZN (n_0_0_264), .A1 (n_0_0_263), .A2 (hfn_ipo_n45), .B1 (n_0_0_235), .B2 (n_0_0_216));
AOI22_X1 i_0_0_352 (.ZN (n_0_0_263), .A1 (n_0_0_262), .A2 (n_0_0_242), .B1 (n_0_0_209), .B2 (n_0_0_244));
NAND2_X1 i_0_0_351 (.ZN (n_0_0_262), .A1 (n_0_0_260), .A2 (n_0_0_261));
AOI22_X1 i_0_0_350 (.ZN (n_0_0_261), .A1 (n_0_0_197), .A2 (\read_data2[11] ), .B1 (\read_data2[10] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_349 (.ZN (n_0_0_260), .A1 (n_0_0_196), .A2 (n_0_14), .B1 (n_0_0_200), .B2 (n_0_44));
OAI22_X1 i_0_0_348 (.ZN (n_0_118), .A1 (n_0_0_253), .A2 (hfn_ipo_n35), .B1 (n_0_0_259), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_347 (.ZN (n_0_0_259), .A1 (n_0_0_258), .A2 (hfn_ipo_n39), .B1 (n_0_0_246), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_346 (.ZN (n_0_0_258), .A1 (n_0_0_257), .A2 (hfn_ipo_n45), .B1 (n_0_0_229), .B2 (n_0_0_216));
AOI22_X1 i_0_0_345 (.ZN (n_0_0_257), .A1 (n_0_0_203), .A2 (n_0_0_244), .B1 (n_0_0_256), .B2 (n_0_0_242));
NAND2_X1 i_0_0_344 (.ZN (n_0_0_256), .A1 (n_0_0_254), .A2 (n_0_0_255));
AOI22_X1 i_0_0_343 (.ZN (n_0_0_255), .A1 (n_0_0_197), .A2 (\read_data2[10] ), .B1 (\read_data2[9] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_342 (.ZN (n_0_0_254), .A1 (n_0_0_196), .A2 (n_0_13), .B1 (n_0_0_200), .B2 (n_0_43));
OAI22_X1 i_0_0_341 (.ZN (n_0_117), .A1 (n_0_0_253), .A2 (hfn_ipo_n49), .B1 (n_0_0_247), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_340 (.ZN (n_0_0_253), .A1 (n_0_0_252), .A2 (hfn_ipo_n39), .B1 (hfn_ipo_n47), .B2 (n_0_0_237));
OAI22_X1 i_0_0_339 (.ZN (n_0_0_252), .A1 (n_0_0_251), .A2 (hfn_ipo_n45), .B1 (n_0_0_222), .B2 (n_0_0_216));
AOI22_X1 i_0_0_338 (.ZN (n_0_0_251), .A1 (n_0_0_242), .A2 (n_0_0_250), .B1 (n_0_0_210), .B2 (n_0_0_244));
NAND2_X1 i_0_0_337 (.ZN (n_0_0_250), .A1 (n_0_0_248), .A2 (n_0_0_249));
AOI22_X1 i_0_0_336 (.ZN (n_0_0_249), .A1 (n_0_0_196), .A2 (n_0_12), .B1 (\read_data2[8] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_335 (.ZN (n_0_0_248), .A1 (n_0_0_197), .A2 (\read_data2[9] ), .B1 (n_0_0_200), .B2 (n_0_42));
OAI22_X1 i_0_0_334 (.ZN (n_0_116), .A1 (n_0_0_238), .A2 (hfn_ipo_n35), .B1 (n_0_0_247), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_333 (.ZN (n_0_0_247), .A1 (n_0_0_246), .A2 (hfn_ipo_n39), .B1 (n_0_0_230), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_332 (.ZN (n_0_0_246), .A1 (n_0_0_245), .A2 (hfn_ipo_n45), .B1 (n_0_0_215), .B2 (n_0_0_216));
AOI22_X1 i_0_0_331 (.ZN (n_0_0_245), .A1 (n_0_0_241), .A2 (n_0_0_242), .B1 (n_0_0_204), .B2 (n_0_0_244));
NOR2_X2 i_0_0_330 (.ZN (n_0_0_244), .A1 (n_0_0_243), .A2 (\shift[4] ));
NAND2_X1 i_0_0_329 (.ZN (n_0_0_243), .A1 (n_0_0_33), .A2 (\shift[3] ));
AND2_X1 i_0_0_328 (.ZN (n_0_0_242), .A1 (n_0_0_172), .A2 (n_0_0_173));
NAND2_X1 i_0_0_327 (.ZN (n_0_0_241), .A1 (n_0_0_239), .A2 (n_0_0_240));
AOI22_X1 i_0_0_326 (.ZN (n_0_0_240), .A1 (n_0_0_196), .A2 (n_0_11), .B1 (\read_data2[7] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_325 (.ZN (n_0_0_239), .A1 (n_0_0_197), .A2 (\read_data2[8] ), .B1 (n_0_0_200), .B2 (n_0_41));
OAI22_X1 i_0_0_324 (.ZN (n_0_115), .A1 (n_0_0_238), .A2 (hfn_ipo_n49), .B1 (n_0_0_231), .B2 (hfn_ipo_n35));
OAI22_X1 i_0_0_323 (.ZN (n_0_0_238), .A1 (n_0_0_223), .A2 (hfn_ipo_n39), .B1 (n_0_0_237), .B2 (hfn_ipo_n47));
OAI22_X1 i_0_0_322 (.ZN (n_0_0_237), .A1 (n_0_0_235), .A2 (n_0_0_174), .B1 (n_0_0_236), .B2 (n_0_0_216));
INV_X1 i_0_0_321 (.ZN (n_0_0_236), .A (n_0_0_209));
INV_X1 i_0_0_320 (.ZN (n_0_0_235), .A (n_0_0_234));
NAND2_X1 i_0_0_319 (.ZN (n_0_0_234), .A1 (n_0_0_232), .A2 (n_0_0_233));
AOI22_X1 i_0_0_318 (.ZN (n_0_0_233), .A1 (n_0_0_196), .A2 (n_0_10), .B1 (\read_data2[6] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_317 (.ZN (n_0_0_232), .A1 (n_0_0_197), .A2 (\read_data2[7] ), .B1 (n_0_0_200), .B2 (n_0_40));
OAI22_X1 i_0_0_316 (.ZN (n_0_114), .A1 (n_0_0_224), .A2 (hfn_ipo_n35), .B1 (n_0_0_231), .B2 (hfn_ipo_n49));
OAI22_X1 i_0_0_315 (.ZN (n_0_0_231), .A1 (n_0_0_230), .A2 (hfn_ipo_n47), .B1 (n_0_0_217), .B2 (hfn_ipo_n39));
OAI22_X1 i_0_0_314 (.ZN (n_0_0_230), .A1 (n_0_0_225), .A2 (n_0_0_216), .B1 (n_0_0_229), .B2 (n_0_0_174));
INV_X1 i_0_0_313 (.ZN (n_0_0_229), .A (n_0_0_228));
NAND2_X1 i_0_0_312 (.ZN (n_0_0_228), .A1 (n_0_0_226), .A2 (n_0_0_227));
AOI22_X1 i_0_0_311 (.ZN (n_0_0_227), .A1 (n_0_0_197), .A2 (\read_data2[6] ), .B1 (\read_data2[5] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_310 (.ZN (n_0_0_226), .A1 (n_0_0_196), .A2 (n_0_9), .B1 (n_0_0_200), .B2 (n_0_39));
INV_X1 i_0_0_309 (.ZN (n_0_0_225), .A (n_0_0_203));
OAI22_X1 i_0_0_308 (.ZN (n_0_113), .A1 (n_0_0_224), .A2 (hfn_ipo_n49), .B1 (n_0_0_218), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_0_307 (.ZN (n_0_0_224), .A1 (n_0_0_223), .A2 (hfn_ipo_n39), .B1 (n_0_0_209), .B2 (n_0_0_205));
OAI22_X1 i_0_0_306 (.ZN (n_0_0_223), .A1 (n_0_0_198), .A2 (n_0_0_216), .B1 (n_0_0_222), .B2 (n_0_0_174));
INV_X1 i_0_0_305 (.ZN (n_0_0_222), .A (n_0_0_221));
NAND2_X1 i_0_0_304 (.ZN (n_0_0_221), .A1 (n_0_0_219), .A2 (n_0_0_220));
AOI22_X1 i_0_0_303 (.ZN (n_0_0_220), .A1 (n_0_0_196), .A2 (n_0_8), .B1 (\read_data2[4] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_302 (.ZN (n_0_0_219), .A1 (n_0_0_197), .A2 (\read_data2[5] ), .B1 (n_0_0_200), .B2 (n_0_38));
OAI22_X1 i_0_0_301 (.ZN (n_0_112), .A1 (n_0_0_218), .A2 (hfn_ipo_n49), .B1 (hfn_ipo_n35), .B2 (n_0_0_211));
AOI22_X1 i_0_0_300 (.ZN (n_0_0_218), .A1 (n_0_0_217), .A2 (hfn_ipo_n39), .B1 (n_0_0_203), .B2 (n_0_0_205));
OAI22_X1 i_0_0_299 (.ZN (n_0_0_217), .A1 (n_0_0_215), .A2 (n_0_0_174), .B1 (n_0_0_171), .B2 (n_0_0_216));
NAND3_X1 i_0_0_298 (.ZN (n_0_0_216), .A1 (n_0_0_172), .A2 (n_0_0_173), .A3 (hfn_ipo_n45));
INV_X1 i_0_0_297 (.ZN (n_0_0_215), .A (n_0_0_214));
NAND2_X1 i_0_0_296 (.ZN (n_0_0_214), .A1 (n_0_0_212), .A2 (n_0_0_213));
AOI22_X1 i_0_0_295 (.ZN (n_0_0_213), .A1 (n_0_0_196), .A2 (n_0_7), .B1 (\read_data2[3] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_294 (.ZN (n_0_0_212), .A1 (n_0_0_197), .A2 (\read_data2[4] ), .B1 (n_0_0_200), .B2 (n_0_37));
AOI22_X1 i_0_0_293 (.ZN (n_0_111), .A1 (n_0_0_211), .A2 (hfn_ipo_n35), .B1 (n_0_0_206), .B2 (hfn_ipo_n49));
AOI22_X1 i_0_0_292 (.ZN (n_0_0_211), .A1 (n_0_0_175), .A2 (n_0_0_209), .B1 (n_0_0_210), .B2 (n_0_0_205));
INV_X1 i_0_0_291 (.ZN (n_0_0_210), .A (n_0_0_198));
NAND2_X1 i_0_0_290 (.ZN (n_0_0_209), .A1 (n_0_0_207), .A2 (n_0_0_208));
AOI22_X1 i_0_0_289 (.ZN (n_0_0_208), .A1 (n_0_0_196), .A2 (n_0_6), .B1 (\read_data2[2] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_288 (.ZN (n_0_0_207), .A1 (n_0_0_197), .A2 (\read_data2[3] ), .B1 (n_0_0_200), .B2 (n_0_36));
OAI22_X2 i_0_0_287 (.ZN (n_0_110), .A1 (n_0_0_198), .A2 (n_0_0_199), .B1 (n_0_0_206), .B2 (hfn_ipo_n49));
AOI22_X2 i_0_0_286 (.ZN (n_0_0_206), .A1 (n_0_0_203), .A2 (n_0_0_175), .B1 (n_0_0_204), .B2 (n_0_0_205));
NOR2_X1 i_0_0_285 (.ZN (n_0_0_205), .A1 (n_0_0_174), .A2 (hfn_ipo_n39));
INV_X1 i_0_0_284 (.ZN (n_0_0_204), .A (n_0_0_171));
NAND2_X2 i_0_0_283 (.ZN (n_0_0_203), .A1 (n_0_0_201), .A2 (n_0_0_202));
AOI22_X2 i_0_0_282 (.ZN (n_0_0_202), .A1 (n_0_0_196), .A2 (n_0_5), .B1 (\read_data2[1] ), .B2 (drc_ipo_n51));
AOI22_X1 i_0_0_281 (.ZN (n_0_0_201), .A1 (n_0_0_197), .A2 (\read_data2[2] ), .B1 (n_0_0_200), .B2 (n_0_35));
INV_X2 i_0_0_280 (.ZN (n_0_0_200), .A (n_0_0_194));
NAND2_X1 i_0_0_279 (.ZN (n_0_0_199), .A1 (n_0_0_175), .A2 (hfn_ipo_n49));
OAI33_X1 i_0_0_278 (.ZN (n_0_109), .A1 (n_0_0_198), .A2 (hfn_ipo_n49), .A3 (n_0_0_176)
    , .B1 (n_0_0_171), .B2 (hfn_ipo_n35), .B3 (n_0_0_176));
AOI221_X2 i_0_0_277 (.ZN (n_0_0_198), .A (n_0_0_195), .B1 (n_0_0_196), .B2 (n_0_4)
    , .C1 (\read_data2[1] ), .C2 (n_0_0_197));
NOR2_X4 i_0_0_276 (.ZN (n_0_0_197), .A1 (n_0_0_169), .A2 (n_0_0_191));
NOR2_X4 i_0_0_275 (.ZN (n_0_0_196), .A1 (n_0_0_169), .A2 (n_0_0_190));
AOI21_X1 i_0_0_274 (.ZN (n_0_0_195), .A (n_0_0_170), .B1 (n_0_0_193), .B2 (n_0_0_194));
NAND3_X1 i_0_0_273 (.ZN (n_0_0_194), .A1 (n_0_0_168), .A2 (n_0_0_166), .A3 (n_0_0_191));
INV_X1 i_0_0_272 (.ZN (n_0_0_193), .A (drc_ipo_n51));
NOR3_X1 i_0_0_271 (.ZN (n_0_0_192), .A1 (n_0_0_168), .A2 (n_0_0_166), .A3 (n_0_0_191));
INV_X1 i_0_0_270 (.ZN (n_0_0_191), .A (n_0_0_190));
AOI211_X1 i_0_0_269 (.ZN (n_0_0_190), .A (n_0_0_183), .B (n_0_0_188), .C1 (n_0_0_123), .C2 (n_0_0_189));
OAI22_X1 i_0_0_268 (.ZN (n_0_0_189), .A1 (n_0_0_120), .A2 (n_0_0_129), .B1 (n_0_0_153), .B2 (n_0_0_138));
AND3_X1 i_0_0_267 (.ZN (n_0_0_188), .A1 (n_0_0_187), .A2 (n_0_0_17), .A3 (\i[2] ));
OAI33_X1 i_0_0_266 (.ZN (n_0_0_187), .A1 (n_0_0_186), .A2 (n_0_0_6), .A3 (n_0_0_1)
    , .B1 (n_0_0_137), .B2 (\i[1] ), .B3 (\i[0] ));
AOI221_X1 i_0_0_265 (.ZN (n_0_0_186), .A (n_0_0_185), .B1 (\read_data[23] ), .B2 (n_0_0_105)
    , .C1 (\read_data[15] ), .C2 (n_0_0_104));
OAI22_X1 i_0_0_264 (.ZN (n_0_0_185), .A1 (n_0_0_160), .A2 (n_0_0_184), .B1 (n_0_0_107), .B2 (n_0_0_118));
INV_X1 i_0_0_263 (.ZN (n_0_0_184), .A (\read_data[7] ));
OAI21_X1 i_0_0_262 (.ZN (n_0_0_183), .A (n_0_0_181), .B1 (n_0_0_130), .B2 (n_0_0_182));
AOI22_X1 i_0_0_261 (.ZN (n_0_0_182), .A1 (n_0_0_110), .A2 (n_0_0_149), .B1 (n_0_0_114), .B2 (n_0_0_144));
AOI221_X1 i_0_0_260 (.ZN (n_0_0_181), .A (n_0_0_178), .B1 (n_0_0_127), .B2 (n_0_0_179)
    , .C1 (n_0_0_180), .C2 (n_0_0_147));
INV_X1 i_0_0_259 (.ZN (n_0_0_180), .A (n_0_0_131));
INV_X1 i_0_0_258 (.ZN (n_0_0_179), .A (n_0_0_124));
NOR3_X1 i_0_0_257 (.ZN (n_0_0_178), .A1 (n_0_0_36), .A2 (\i[5] ), .A3 (n_0_0_177));
INV_X1 i_0_0_256 (.ZN (n_0_0_177), .A (\read_data[0] ));
NOR3_X1 i_0_0_255 (.ZN (n_0_108), .A1 (n_0_0_171), .A2 (hfn_ipo_n49), .A3 (n_0_0_176));
INV_X1 i_0_0_254 (.ZN (n_0_0_176), .A (n_0_0_175));
NOR2_X1 i_0_0_253 (.ZN (n_0_0_175), .A1 (n_0_0_174), .A2 (hfn_ipo_n47));
NAND3_X1 i_0_0_252 (.ZN (n_0_0_174), .A1 (n_0_0_172), .A2 (n_0_0_173), .A3 (hfn_ipo_n37));
INV_X1 i_0_0_251 (.ZN (n_0_0_173), .A (\shift[4] ));
NOR2_X2 i_0_0_250 (.ZN (n_0_0_172), .A1 (\shift[5] ), .A2 (\shift[3] ));
OR2_X1 i_0_0_249 (.ZN (n_0_0_171), .A1 (n_0_0_169), .A2 (n_0_0_170));
INV_X1 i_0_0_248 (.ZN (n_0_0_170), .A (\read_data2[0] ));
OAI22_X2 i_0_0_247 (.ZN (n_0_0_169), .A1 (n_0_0_151), .A2 (n_0_0_167), .B1 (n_0_0_168), .B2 (n_0_0_166));
INV_X1 i_0_0_246 (.ZN (n_0_0_168), .A (n_0_0_151));
INV_X1 i_0_0_245 (.ZN (n_0_0_167), .A (n_0_0_166));
NOR2_X1 i_0_0_244 (.ZN (n_0_0_166), .A1 (n_0_0_164), .A2 (n_0_0_165));
OAI22_X1 i_0_0_243 (.ZN (n_0_0_165), .A1 (n_0_0_122), .A2 (n_0_0_131), .B1 (n_0_0_124), .B2 (n_0_0_133));
OAI211_X1 i_0_0_242 (.ZN (n_0_0_164), .A (n_0_0_155), .B (n_0_0_162), .C1 (n_0_0_130), .C2 (n_0_0_163));
AOI22_X1 i_0_0_241 (.ZN (n_0_0_163), .A1 (n_0_0_127), .A2 (n_0_0_149), .B1 (n_0_0_136), .B2 (n_0_0_144));
AOI22_X1 i_0_0_240 (.ZN (n_0_0_162), .A1 (n_0_0_157), .A2 (n_0_0_123), .B1 (n_0_0_159), .B2 (n_0_0_161));
NOR3_X1 i_0_0_239 (.ZN (n_0_0_161), .A1 (n_0_0_160), .A2 (n_0_0_17), .A3 (\i[1] ));
INV_X1 i_0_0_238 (.ZN (n_0_0_160), .A (n_0_0_35));
OAI22_X1 i_0_0_237 (.ZN (n_0_0_159), .A1 (n_0_0_129), .A2 (n_0_0_158), .B1 (n_0_0_148), .B2 (n_0_0_118));
INV_X1 i_0_0_236 (.ZN (n_0_0_158), .A (\read_data[30] ));
OAI22_X1 i_0_0_235 (.ZN (n_0_0_157), .A1 (n_0_0_156), .A2 (n_0_0_129), .B1 (n_0_0_111), .B2 (n_0_0_138));
AOI222_X1 i_0_0_234 (.ZN (n_0_0_156), .A1 (\read_data[22] ), .A2 (n_0_0_108), .B1 (n_0_0_105)
    , .B2 (\read_data[14] ), .C1 (n_0_0_104), .C2 (\read_data[6] ));
NAND3_X1 i_0_0_233 (.ZN (n_0_0_155), .A1 (n_0_0_154), .A2 (n_0_0_17), .A3 (\i[2] ));
OAI33_X1 i_0_0_232 (.ZN (n_0_0_154), .A1 (n_0_0_152), .A2 (\i[1] ), .A3 (\i[0] ), .B1 (n_0_0_153)
    , .B2 (n_0_0_6), .B3 (n_0_0_1));
INV_X1 i_0_0_231 (.ZN (n_0_0_153), .A (n_0_0_143));
INV_X1 i_0_0_230 (.ZN (n_0_0_152), .A (n_0_0_147));
OAI211_X1 i_0_0_229 (.ZN (n_0_0_151), .A (n_0_0_117), .B (n_0_0_140), .C1 (n_0_0_130), .C2 (n_0_0_150));
AOI22_X1 i_0_0_228 (.ZN (n_0_0_150), .A1 (n_0_0_143), .A2 (n_0_0_144), .B1 (n_0_0_147), .B2 (n_0_0_149));
INV_X1 i_0_0_227 (.ZN (n_0_0_149), .A (n_0_0_148));
NAND2_X1 i_0_0_226 (.ZN (n_0_0_148), .A1 (n_0_0_7), .A2 (\i[0] ));
NAND2_X1 i_0_0_225 (.ZN (n_0_0_147), .A1 (n_0_0_145), .A2 (n_0_0_146));
AOI22_X1 i_0_0_224 (.ZN (n_0_0_146), .A1 (n_0_0_108), .A2 (\read_data[26] ), .B1 (n_0_0_35), .B2 (\read_data[2] ));
AOI22_X1 i_0_0_223 (.ZN (n_0_0_145), .A1 (n_0_0_104), .A2 (\read_data[10] ), .B1 (n_0_0_105), .B2 (\read_data[18] ));
NOR2_X1 i_0_0_222 (.ZN (n_0_0_144), .A1 (n_0_0_7), .A2 (\i[0] ));
NAND2_X1 i_0_0_221 (.ZN (n_0_0_143), .A1 (n_0_0_141), .A2 (n_0_0_142));
AOI22_X1 i_0_0_220 (.ZN (n_0_0_142), .A1 (n_0_0_108), .A2 (\read_data[29] ), .B1 (n_0_0_35), .B2 (\read_data[5] ));
AOI22_X1 i_0_0_219 (.ZN (n_0_0_141), .A1 (n_0_0_104), .A2 (\read_data[13] ), .B1 (n_0_0_105), .B2 (\read_data[21] ));
AOI211_X1 i_0_0_218 (.ZN (n_0_0_140), .A (n_0_0_119), .B (n_0_0_132), .C1 (n_0_0_123), .C2 (n_0_0_139));
OAI22_X1 i_0_0_217 (.ZN (n_0_0_139), .A1 (n_0_0_133), .A2 (n_0_0_129), .B1 (n_0_0_137), .B2 (n_0_0_138));
NAND2_X1 i_0_0_216 (.ZN (n_0_0_138), .A1 (\i[0] ), .A2 (\i[2] ));
INV_X1 i_0_0_215 (.ZN (n_0_0_137), .A (n_0_0_136));
NAND2_X1 i_0_0_214 (.ZN (n_0_0_136), .A1 (n_0_0_134), .A2 (n_0_0_135));
AOI22_X1 i_0_0_213 (.ZN (n_0_0_135), .A1 (n_0_0_108), .A2 (\read_data[28] ), .B1 (n_0_0_35), .B2 (\read_data[4] ));
AOI22_X1 i_0_0_212 (.ZN (n_0_0_134), .A1 (n_0_0_104), .A2 (\read_data[12] ), .B1 (n_0_0_105), .B2 (\read_data[20] ));
AOI222_X1 i_0_0_211 (.ZN (n_0_0_133), .A1 (n_0_0_108), .A2 (\read_data[23] ), .B1 (n_0_0_105)
    , .B2 (\read_data[15] ), .C1 (n_0_0_104), .C2 (\read_data[7] ));
OAI22_X1 i_0_0_210 (.ZN (n_0_0_132), .A1 (n_0_0_122), .A2 (n_0_0_124), .B1 (n_0_0_128), .B2 (n_0_0_131));
OR2_X1 i_0_0_209 (.ZN (n_0_0_131), .A1 (n_0_0_129), .A2 (n_0_0_130));
NAND2_X1 i_0_0_208 (.ZN (n_0_0_130), .A1 (n_0_0_17), .A2 (\i[1] ));
INV_X1 i_0_0_207 (.ZN (n_0_0_129), .A (n_0_0_34));
INV_X1 i_0_0_206 (.ZN (n_0_0_128), .A (n_0_0_127));
NAND2_X1 i_0_0_205 (.ZN (n_0_0_127), .A1 (n_0_0_125), .A2 (n_0_0_126));
AOI22_X1 i_0_0_204 (.ZN (n_0_0_126), .A1 (n_0_0_108), .A2 (\read_data[25] ), .B1 (n_0_0_35), .B2 (\read_data[1] ));
AOI22_X1 i_0_0_203 (.ZN (n_0_0_125), .A1 (n_0_0_104), .A2 (\read_data[9] ), .B1 (n_0_0_105), .B2 (\read_data[17] ));
NAND3_X1 i_0_0_202 (.ZN (n_0_0_124), .A1 (n_0_0_123), .A2 (\i[0] ), .A3 (n_0_0_7));
NOR2_X1 i_0_0_201 (.ZN (n_0_0_123), .A1 (\i[5] ), .A2 (\i[1] ));
AOI21_X1 i_0_0_200 (.ZN (n_0_0_122), .A (n_0_0_121), .B1 (\read_data[0] ), .B2 (n_0_0_35));
INV_X1 i_0_0_199 (.ZN (n_0_0_121), .A (n_0_0_120));
AOI222_X1 i_0_0_198 (.ZN (n_0_0_120), .A1 (n_0_0_108), .A2 (\read_data[24] ), .B1 (n_0_0_104)
    , .B2 (\read_data[8] ), .C1 (n_0_0_105), .C2 (\read_data[16] ));
NOR3_X1 i_0_0_197 (.ZN (n_0_0_119), .A1 (n_0_0_36), .A2 (n_0_0_17), .A3 (n_0_0_118));
INV_X1 i_0_0_196 (.ZN (n_0_0_118), .A (\read_data[31] ));
NAND3_X1 i_0_0_195 (.ZN (n_0_0_117), .A1 (n_0_0_116), .A2 (n_0_0_17), .A3 (\i[2] ));
OAI33_X1 i_0_0_194 (.ZN (n_0_0_116), .A1 (n_0_0_111), .A2 (\i[1] ), .A3 (\i[0] ), .B1 (n_0_0_115)
    , .B2 (n_0_0_6), .B3 (n_0_0_1));
INV_X1 i_0_0_193 (.ZN (n_0_0_115), .A (n_0_0_114));
NAND2_X1 i_0_0_192 (.ZN (n_0_0_114), .A1 (n_0_0_112), .A2 (n_0_0_113));
AOI22_X1 i_0_0_191 (.ZN (n_0_0_113), .A1 (n_0_0_108), .A2 (\read_data[30] ), .B1 (n_0_0_35), .B2 (\read_data[6] ));
AOI22_X1 i_0_0_190 (.ZN (n_0_0_112), .A1 (n_0_0_104), .A2 (\read_data[14] ), .B1 (n_0_0_105), .B2 (\read_data[22] ));
INV_X1 i_0_0_189 (.ZN (n_0_0_111), .A (n_0_0_110));
NAND2_X1 i_0_0_188 (.ZN (n_0_0_110), .A1 (n_0_0_106), .A2 (n_0_0_109));
AOI22_X1 i_0_0_187 (.ZN (n_0_0_109), .A1 (n_0_0_108), .A2 (\read_data[27] ), .B1 (n_0_0_35), .B2 (\read_data[3] ));
INV_X2 i_0_0_186 (.ZN (n_0_0_108), .A (n_0_0_107));
NAND2_X1 i_0_0_185 (.ZN (n_0_0_107), .A1 (\i[4] ), .A2 (\i[3] ));
AOI22_X1 i_0_0_184 (.ZN (n_0_0_106), .A1 (n_0_0_104), .A2 (\read_data[11] ), .B1 (n_0_0_105), .B2 (\read_data[19] ));
NOR2_X2 i_0_0_183 (.ZN (n_0_0_105), .A1 (n_0_0_103), .A2 (\i[3] ));
AND2_X2 i_0_0_182 (.ZN (n_0_0_104), .A1 (n_0_0_103), .A2 (\i[3] ));
INV_X2 i_0_0_181 (.ZN (n_0_0_103), .A (\i[4] ));
INV_X1 i_0_0_180 (.ZN (n_0_104), .A (n_0_0_102));
AOI22_X1 i_0_0_179 (.ZN (n_0_0_102), .A1 (hfn_ipo_n41), .A2 (n_0_234), .B1 (hfn_ipo_n43), .B2 (\res[63] ));
INV_X1 i_0_0_178 (.ZN (n_0_103), .A (n_0_0_101));
AOI22_X1 i_0_0_177 (.ZN (n_0_0_101), .A1 (hfn_ipo_n41), .A2 (n_0_233), .B1 (hfn_ipo_n43), .B2 (\res[62] ));
INV_X1 i_0_0_176 (.ZN (n_0_102), .A (n_0_0_100));
AOI22_X1 i_0_0_175 (.ZN (n_0_0_100), .A1 (hfn_ipo_n41), .A2 (n_0_232), .B1 (hfn_ipo_n43), .B2 (\res[61] ));
INV_X1 i_0_0_174 (.ZN (n_0_101), .A (n_0_0_99));
AOI22_X1 i_0_0_173 (.ZN (n_0_0_99), .A1 (hfn_ipo_n41), .A2 (n_0_231), .B1 (hfn_ipo_n43), .B2 (\res[60] ));
INV_X1 i_0_0_172 (.ZN (n_0_100), .A (n_0_0_98));
AOI22_X1 i_0_0_171 (.ZN (n_0_0_98), .A1 (hfn_ipo_n41), .A2 (n_0_230), .B1 (hfn_ipo_n43), .B2 (\res[59] ));
INV_X1 i_0_0_170 (.ZN (n_0_99), .A (n_0_0_97));
AOI22_X1 i_0_0_169 (.ZN (n_0_0_97), .A1 (hfn_ipo_n41), .A2 (n_0_229), .B1 (hfn_ipo_n43), .B2 (\res[58] ));
INV_X1 i_0_0_168 (.ZN (n_0_98), .A (n_0_0_96));
AOI22_X1 i_0_0_167 (.ZN (n_0_0_96), .A1 (hfn_ipo_n41), .A2 (n_0_228), .B1 (hfn_ipo_n43), .B2 (\res[57] ));
INV_X1 i_0_0_166 (.ZN (n_0_97), .A (n_0_0_95));
AOI22_X1 i_0_0_165 (.ZN (n_0_0_95), .A1 (hfn_ipo_n41), .A2 (n_0_227), .B1 (hfn_ipo_n43), .B2 (\res[56] ));
INV_X1 i_0_0_164 (.ZN (n_0_96), .A (n_0_0_94));
AOI22_X1 i_0_0_163 (.ZN (n_0_0_94), .A1 (hfn_ipo_n41), .A2 (n_0_226), .B1 (hfn_ipo_n43), .B2 (\res[55] ));
INV_X1 i_0_0_162 (.ZN (n_0_95), .A (n_0_0_93));
AOI22_X1 i_0_0_161 (.ZN (n_0_0_93), .A1 (hfn_ipo_n41), .A2 (n_0_225), .B1 (hfn_ipo_n43), .B2 (\res[54] ));
INV_X1 i_0_0_160 (.ZN (n_0_94), .A (n_0_0_92));
AOI22_X1 i_0_0_159 (.ZN (n_0_0_92), .A1 (hfn_ipo_n41), .A2 (n_0_224), .B1 (hfn_ipo_n43), .B2 (\res[53] ));
INV_X1 i_0_0_158 (.ZN (n_0_93), .A (n_0_0_91));
AOI22_X1 i_0_0_157 (.ZN (n_0_0_91), .A1 (hfn_ipo_n41), .A2 (n_0_223), .B1 (hfn_ipo_n43), .B2 (\res[52] ));
INV_X1 i_0_0_156 (.ZN (n_0_92), .A (n_0_0_90));
AOI22_X1 i_0_0_155 (.ZN (n_0_0_90), .A1 (hfn_ipo_n41), .A2 (n_0_222), .B1 (hfn_ipo_n43), .B2 (\res[51] ));
INV_X1 i_0_0_154 (.ZN (n_0_91), .A (n_0_0_89));
AOI22_X1 i_0_0_153 (.ZN (n_0_0_89), .A1 (hfn_ipo_n41), .A2 (n_0_221), .B1 (hfn_ipo_n43), .B2 (\res[50] ));
INV_X1 i_0_0_152 (.ZN (n_0_90), .A (n_0_0_88));
AOI22_X1 i_0_0_151 (.ZN (n_0_0_88), .A1 (hfn_ipo_n41), .A2 (n_0_220), .B1 (hfn_ipo_n43), .B2 (\res[49] ));
INV_X1 i_0_0_150 (.ZN (n_0_89), .A (n_0_0_87));
AOI22_X1 i_0_0_149 (.ZN (n_0_0_87), .A1 (n_0_105), .A2 (n_0_219), .B1 (hfn_ipo_n44), .B2 (\res[48] ));
INV_X1 i_0_0_148 (.ZN (n_0_88), .A (n_0_0_86));
AOI22_X1 i_0_0_147 (.ZN (n_0_0_86), .A1 (n_0_105), .A2 (n_0_218), .B1 (hfn_ipo_n44), .B2 (\res[47] ));
INV_X1 i_0_0_146 (.ZN (n_0_87), .A (n_0_0_85));
AOI22_X1 i_0_0_145 (.ZN (n_0_0_85), .A1 (n_0_105), .A2 (n_0_217), .B1 (hfn_ipo_n44), .B2 (\res[46] ));
INV_X1 i_0_0_144 (.ZN (n_0_86), .A (n_0_0_84));
AOI22_X1 i_0_0_143 (.ZN (n_0_0_84), .A1 (n_0_105), .A2 (n_0_216), .B1 (hfn_ipo_n44), .B2 (\res[45] ));
INV_X1 i_0_0_142 (.ZN (n_0_85), .A (n_0_0_83));
AOI22_X1 i_0_0_141 (.ZN (n_0_0_83), .A1 (n_0_105), .A2 (n_0_215), .B1 (hfn_ipo_n44), .B2 (\res[44] ));
INV_X1 i_0_0_140 (.ZN (n_0_84), .A (n_0_0_82));
AOI22_X1 i_0_0_139 (.ZN (n_0_0_82), .A1 (n_0_105), .A2 (n_0_214), .B1 (hfn_ipo_n44), .B2 (\res[43] ));
INV_X1 i_0_0_138 (.ZN (n_0_83), .A (n_0_0_81));
AOI22_X1 i_0_0_137 (.ZN (n_0_0_81), .A1 (n_0_105), .A2 (n_0_213), .B1 (hfn_ipo_n44), .B2 (\res[42] ));
INV_X1 i_0_0_136 (.ZN (n_0_82), .A (n_0_0_80));
AOI22_X1 i_0_0_135 (.ZN (n_0_0_80), .A1 (n_0_105), .A2 (n_0_212), .B1 (hfn_ipo_n44), .B2 (\res[41] ));
INV_X1 i_0_0_134 (.ZN (n_0_81), .A (n_0_0_79));
AOI22_X1 i_0_0_133 (.ZN (n_0_0_79), .A1 (n_0_105), .A2 (n_0_211), .B1 (hfn_ipo_n44), .B2 (\res[40] ));
INV_X1 i_0_0_132 (.ZN (n_0_80), .A (n_0_0_78));
AOI22_X1 i_0_0_131 (.ZN (n_0_0_78), .A1 (n_0_105), .A2 (n_0_210), .B1 (hfn_ipo_n44), .B2 (\res[39] ));
INV_X1 i_0_0_130 (.ZN (n_0_79), .A (n_0_0_77));
AOI22_X1 i_0_0_129 (.ZN (n_0_0_77), .A1 (n_0_105), .A2 (n_0_209), .B1 (hfn_ipo_n44), .B2 (\res[38] ));
INV_X1 i_0_0_128 (.ZN (n_0_78), .A (n_0_0_76));
AOI22_X1 i_0_0_127 (.ZN (n_0_0_76), .A1 (n_0_105), .A2 (n_0_208), .B1 (hfn_ipo_n44), .B2 (\res[37] ));
INV_X1 i_0_0_126 (.ZN (n_0_77), .A (n_0_0_75));
AOI22_X1 i_0_0_125 (.ZN (n_0_0_75), .A1 (n_0_105), .A2 (n_0_207), .B1 (hfn_ipo_n44), .B2 (\res[36] ));
INV_X1 i_0_0_124 (.ZN (n_0_76), .A (n_0_0_74));
AOI22_X1 i_0_0_123 (.ZN (n_0_0_74), .A1 (n_0_105), .A2 (n_0_206), .B1 (hfn_ipo_n44), .B2 (\res[35] ));
INV_X1 i_0_0_122 (.ZN (n_0_269), .A (n_0_0_73));
AOI22_X1 i_0_0_121 (.ZN (n_0_0_73), .A1 (n_0_105), .A2 (n_0_205), .B1 (hfn_ipo_n44), .B2 (\res[34] ));
INV_X1 i_0_0_120 (.ZN (n_0_268), .A (n_0_0_72));
AOI22_X1 i_0_0_119 (.ZN (n_0_0_72), .A1 (n_0_105), .A2 (n_0_204), .B1 (hfn_ipo_n44), .B2 (\res[33] ));
INV_X1 i_0_0_118 (.ZN (n_0_267), .A (n_0_0_71));
AOI22_X1 i_0_0_117 (.ZN (n_0_0_71), .A1 (n_0_105), .A2 (n_0_203), .B1 (hfn_ipo_n44), .B2 (\res[32] ));
INV_X1 i_0_0_116 (.ZN (n_0_266), .A (n_0_0_70));
AOI22_X1 i_0_0_115 (.ZN (n_0_0_70), .A1 (n_0_105), .A2 (n_0_202), .B1 (hfn_ipo_n44), .B2 (\res[31] ));
INV_X1 i_0_0_114 (.ZN (n_0_265), .A (n_0_0_69));
AOI22_X1 i_0_0_113 (.ZN (n_0_0_69), .A1 (n_0_105), .A2 (n_0_201), .B1 (hfn_ipo_n44), .B2 (\res[30] ));
INV_X1 i_0_0_112 (.ZN (n_0_264), .A (n_0_0_68));
AOI22_X1 i_0_0_111 (.ZN (n_0_0_68), .A1 (n_0_105), .A2 (n_0_200), .B1 (hfn_ipo_n44), .B2 (\res[29] ));
INV_X1 i_0_0_110 (.ZN (n_0_263), .A (n_0_0_67));
AOI22_X1 i_0_0_109 (.ZN (n_0_0_67), .A1 (n_0_105), .A2 (n_0_199), .B1 (hfn_ipo_n44), .B2 (\res[28] ));
INV_X1 i_0_0_108 (.ZN (n_0_262), .A (n_0_0_66));
AOI22_X1 i_0_0_107 (.ZN (n_0_0_66), .A1 (n_0_105), .A2 (n_0_198), .B1 (hfn_ipo_n44), .B2 (\res[27] ));
INV_X1 i_0_0_106 (.ZN (n_0_261), .A (n_0_0_65));
AOI22_X1 i_0_0_105 (.ZN (n_0_0_65), .A1 (n_0_105), .A2 (n_0_197), .B1 (hfn_ipo_n44), .B2 (\res[26] ));
INV_X1 i_0_0_104 (.ZN (n_0_260), .A (n_0_0_64));
AOI22_X1 i_0_0_103 (.ZN (n_0_0_64), .A1 (hfn_ipo_n41), .A2 (n_0_196), .B1 (hfn_ipo_n43), .B2 (\res[25] ));
INV_X1 i_0_0_102 (.ZN (n_0_259), .A (n_0_0_63));
AOI22_X1 i_0_0_101 (.ZN (n_0_0_63), .A1 (hfn_ipo_n41), .A2 (n_0_195), .B1 (hfn_ipo_n43), .B2 (\res[24] ));
INV_X1 i_0_0_100 (.ZN (n_0_258), .A (n_0_0_62));
AOI22_X1 i_0_0_99 (.ZN (n_0_0_62), .A1 (hfn_ipo_n41), .A2 (n_0_194), .B1 (hfn_ipo_n43), .B2 (\res[23] ));
INV_X1 i_0_0_98 (.ZN (n_0_257), .A (n_0_0_61));
AOI22_X1 i_0_0_97 (.ZN (n_0_0_61), .A1 (hfn_ipo_n41), .A2 (n_0_193), .B1 (hfn_ipo_n43), .B2 (\res[22] ));
INV_X1 i_0_0_96 (.ZN (n_0_256), .A (n_0_0_60));
AOI22_X1 i_0_0_95 (.ZN (n_0_0_60), .A1 (hfn_ipo_n41), .A2 (n_0_192), .B1 (hfn_ipo_n43), .B2 (\res[21] ));
INV_X1 i_0_0_94 (.ZN (n_0_255), .A (n_0_0_59));
AOI22_X1 i_0_0_93 (.ZN (n_0_0_59), .A1 (hfn_ipo_n41), .A2 (n_0_191), .B1 (hfn_ipo_n43), .B2 (\res[20] ));
INV_X1 i_0_0_92 (.ZN (n_0_254), .A (n_0_0_58));
AOI22_X1 i_0_0_91 (.ZN (n_0_0_58), .A1 (hfn_ipo_n41), .A2 (n_0_190), .B1 (hfn_ipo_n43), .B2 (\res[19] ));
INV_X1 i_0_0_90 (.ZN (n_0_253), .A (n_0_0_57));
AOI22_X1 i_0_0_89 (.ZN (n_0_0_57), .A1 (hfn_ipo_n41), .A2 (n_0_189), .B1 (hfn_ipo_n43), .B2 (\res[18] ));
INV_X1 i_0_0_88 (.ZN (n_0_252), .A (n_0_0_56));
AOI22_X1 i_0_0_87 (.ZN (n_0_0_56), .A1 (hfn_ipo_n41), .A2 (n_0_188), .B1 (hfn_ipo_n43), .B2 (\res[17] ));
INV_X1 i_0_0_86 (.ZN (n_0_251), .A (n_0_0_55));
AOI22_X1 i_0_0_85 (.ZN (n_0_0_55), .A1 (hfn_ipo_n41), .A2 (n_0_187), .B1 (hfn_ipo_n43), .B2 (\res[16] ));
INV_X1 i_0_0_84 (.ZN (n_0_250), .A (n_0_0_54));
AOI22_X1 i_0_0_83 (.ZN (n_0_0_54), .A1 (hfn_ipo_n41), .A2 (n_0_186), .B1 (hfn_ipo_n43), .B2 (\res[15] ));
INV_X1 i_0_0_82 (.ZN (n_0_249), .A (n_0_0_53));
AOI22_X1 i_0_0_81 (.ZN (n_0_0_53), .A1 (hfn_ipo_n41), .A2 (n_0_185), .B1 (hfn_ipo_n43), .B2 (\res[14] ));
INV_X1 i_0_0_80 (.ZN (n_0_248), .A (n_0_0_52));
AOI22_X1 i_0_0_79 (.ZN (n_0_0_52), .A1 (hfn_ipo_n41), .A2 (n_0_184), .B1 (hfn_ipo_n43), .B2 (\res[13] ));
INV_X1 i_0_0_78 (.ZN (n_0_247), .A (n_0_0_51));
AOI22_X1 i_0_0_77 (.ZN (n_0_0_51), .A1 (hfn_ipo_n41), .A2 (n_0_183), .B1 (hfn_ipo_n43), .B2 (\res[12] ));
INV_X1 i_0_0_76 (.ZN (n_0_246), .A (n_0_0_50));
AOI22_X1 i_0_0_75 (.ZN (n_0_0_50), .A1 (hfn_ipo_n41), .A2 (n_0_182), .B1 (hfn_ipo_n43), .B2 (\res[11] ));
INV_X1 i_0_0_74 (.ZN (n_0_245), .A (n_0_0_49));
AOI22_X1 i_0_0_73 (.ZN (n_0_0_49), .A1 (hfn_ipo_n41), .A2 (n_0_181), .B1 (hfn_ipo_n43), .B2 (\res[10] ));
INV_X1 i_0_0_72 (.ZN (n_0_244), .A (n_0_0_48));
AOI22_X1 i_0_0_71 (.ZN (n_0_0_48), .A1 (hfn_ipo_n41), .A2 (n_0_180), .B1 (hfn_ipo_n43), .B2 (\res[9] ));
INV_X1 i_0_0_70 (.ZN (n_0_243), .A (n_0_0_47));
AOI22_X1 i_0_0_69 (.ZN (n_0_0_47), .A1 (hfn_ipo_n41), .A2 (n_0_179), .B1 (hfn_ipo_n43), .B2 (\res[8] ));
INV_X1 i_0_0_68 (.ZN (n_0_242), .A (n_0_0_46));
AOI22_X1 i_0_0_67 (.ZN (n_0_0_46), .A1 (hfn_ipo_n41), .A2 (n_0_178), .B1 (hfn_ipo_n43), .B2 (\res[7] ));
INV_X1 i_0_0_66 (.ZN (n_0_241), .A (n_0_0_45));
AOI22_X1 i_0_0_65 (.ZN (n_0_0_45), .A1 (hfn_ipo_n41), .A2 (n_0_177), .B1 (hfn_ipo_n43), .B2 (\res[6] ));
INV_X1 i_0_0_64 (.ZN (n_0_240), .A (n_0_0_44));
AOI22_X1 i_0_0_63 (.ZN (n_0_0_44), .A1 (hfn_ipo_n41), .A2 (n_0_176), .B1 (hfn_ipo_n43), .B2 (\res[5] ));
INV_X1 i_0_0_62 (.ZN (n_0_239), .A (n_0_0_43));
AOI22_X1 i_0_0_61 (.ZN (n_0_0_43), .A1 (hfn_ipo_n41), .A2 (n_0_175), .B1 (hfn_ipo_n43), .B2 (\res[4] ));
INV_X1 i_0_0_60 (.ZN (n_0_238), .A (n_0_0_42));
AOI22_X1 i_0_0_59 (.ZN (n_0_0_42), .A1 (hfn_ipo_n41), .A2 (n_0_174), .B1 (hfn_ipo_n43), .B2 (\res[3] ));
INV_X1 i_0_0_58 (.ZN (n_0_237), .A (n_0_0_41));
AOI22_X1 i_0_0_57 (.ZN (n_0_0_41), .A1 (hfn_ipo_n41), .A2 (n_0_173), .B1 (hfn_ipo_n43), .B2 (\res[2] ));
INV_X1 i_0_0_56 (.ZN (n_0_236), .A (n_0_0_40));
AOI22_X1 i_0_0_55 (.ZN (n_0_0_40), .A1 (hfn_ipo_n41), .A2 (n_0_172), .B1 (hfn_ipo_n43), .B2 (\res[1] ));
INV_X1 i_0_0_54 (.ZN (n_0_235), .A (n_0_0_39));
AOI22_X1 i_0_0_53 (.ZN (n_0_0_39), .A1 (hfn_ipo_n41), .A2 (n_0_171), .B1 (hfn_ipo_n43), .B2 (\res[0] ));
INV_X1 i_0_0_52 (.ZN (n_0_69), .A (hfn_ipo_n43));
NOR2_X1 i_0_0_51 (.ZN (n_0_0_38), .A1 (n_0_0_37), .A2 (CLOCK_slh_n298));
AND2_X1 i_0_0_50 (.ZN (n_0_105), .A1 (n_0_0_37), .A2 (n_0_0_4));
NAND2_X1 i_0_0_49 (.ZN (n_0_0_37), .A1 (n_0_0_36), .A2 (\i[5] ));
NAND3_X1 i_0_0_48 (.ZN (n_0_0_36), .A1 (n_0_0_34), .A2 (n_0_0_35), .A3 (n_0_0_6));
NOR2_X2 i_0_0_47 (.ZN (n_0_0_35), .A1 (\i[4] ), .A2 (\i[3] ));
NOR2_X1 i_0_0_46 (.ZN (n_0_0_34), .A1 (\i[0] ), .A2 (\i[2] ));
AOI221_X1 i_0_0_45 (.ZN (n_0_75), .A (CLOCK_slh_n298), .B1 (n_0_0_32), .B2 (\shift[5] )
    , .C1 (n_0_0_33), .C2 (n_0_0_31));
INV_X1 i_0_0_44 (.ZN (n_0_0_33), .A (\shift[5] ));
OAI21_X1 i_0_0_43 (.ZN (CLOCK_slh__n635), .A (n_0_0_29), .B1 (n_0_0_30), .B2 (n_0_0_32));
INV_X1 i_0_0_42 (.ZN (n_0_0_32), .A (n_0_0_31));
NAND2_X1 i_0_0_41 (.ZN (n_0_0_31), .A1 (n_0_0_28), .A2 (\shift[4] ));
OAI21_X1 i_0_0_40 (.ZN (n_0_0_30), .A (n_0_0_4), .B1 (n_0_0_28), .B2 (\shift[4] ));
NAND2_X1 i_0_0_39 (.ZN (n_0_0_29), .A1 (start_shift[4]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_38 (.ZN (CLOCK_slh__n633), .A (n_0_0_26), .B1 (n_0_0_27), .B2 (n_0_0_28));
AND2_X1 i_0_0_37 (.ZN (n_0_0_28), .A1 (n_0_0_25), .A2 (\shift[3] ));
OAI21_X1 i_0_0_36 (.ZN (n_0_0_27), .A (n_0_0_4), .B1 (n_0_0_25), .B2 (\shift[3] ));
NAND2_X1 i_0_0_35 (.ZN (n_0_0_26), .A1 (start_shift[3]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_34 (.ZN (CLOCK_slh__n637), .A (n_0_0_21), .B1 (n_0_0_22), .B2 (n_0_0_25));
NOR2_X1 i_0_0_33 (.ZN (n_0_0_25), .A1 (hfn_ipo_n37), .A2 (hfn_ipo_n39));
INV_X1 i_0_0_32 (.ZN (n_0_0_24), .A (hfn_ipo_n47));
INV_X1 i_0_0_31 (.ZN (n_0_0_23), .A (hfn_ipo_n45));
OAI21_X1 i_0_0_30 (.ZN (n_0_0_22), .A (n_0_0_4), .B1 (hfn_ipo_n45), .B2 (hfn_ipo_n47));
NAND2_X1 i_0_0_29 (.ZN (n_0_0_21), .A1 (start_shift[2]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_28 (.ZN (CLOCK_slh__n619), .A (n_0_0_20), .B1 (CLOCK_slh_n298), .B2 (hfn_ipo_n47));
NAND2_X1 i_0_0_27 (.ZN (n_0_0_20), .A1 (start_shift[1]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_26 (.ZN (CLOCK_slh__n625), .A (n_0_0_18), .B1 (hfn_ipo_n35), .B2 (CLOCK_slh_n298));
INV_X1 i_0_0_25 (.ZN (n_0_0_19), .A (hfn_ipo_n49));
NAND2_X1 i_0_0_24 (.ZN (n_0_0_18), .A1 (start_shift[0]), .A2 (CLOCK_slh_n298));
AOI221_X1 i_0_0_23 (.ZN (n_0_68), .A (CLOCK_slh_n298), .B1 (n_0_0_16), .B2 (\i[5] )
    , .C1 (n_0_0_17), .C2 (n_0_0_15));
INV_X1 i_0_0_22 (.ZN (n_0_0_17), .A (\i[5] ));
OAI21_X1 i_0_0_21 (.ZN (CLOCK_slh__n631), .A (n_0_0_12), .B1 (n_0_0_14), .B2 (n_0_0_16));
INV_X1 i_0_0_20 (.ZN (n_0_0_16), .A (n_0_0_15));
NAND2_X1 i_0_0_19 (.ZN (n_0_0_15), .A1 (n_0_0_13), .A2 (\i[4] ));
OAI21_X1 i_0_0_18 (.ZN (n_0_0_14), .A (n_0_0_4), .B1 (n_0_0_13), .B2 (\i[4] ));
INV_X1 i_0_0_17 (.ZN (n_0_0_13), .A (n_0_0_9));
NAND2_X1 i_0_0_16 (.ZN (n_0_0_12), .A1 (start_i[4]), .A2 (CLOCK_slh_n298));
AOI22_X1 i_0_0_15 (.ZN (CLOCK_slh__n627), .A1 (n_0_0_10), .A2 (n_0_0_4), .B1 (n_0_0_11), .B2 (CLOCK_slh_n298));
INV_X1 i_0_0_14 (.ZN (n_0_0_11), .A (start_i[3]));
OAI21_X1 i_0_0_13 (.ZN (n_0_0_10), .A (n_0_0_9), .B1 (\i[3] ), .B2 (n_0_0_8));
NAND2_X1 i_0_0_12 (.ZN (n_0_0_9), .A1 (n_0_0_8), .A2 (\i[3] ));
OAI21_X1 i_0_0_11 (.ZN (CLOCK_slh__n629), .A (n_0_0_3), .B1 (n_0_0_5), .B2 (n_0_0_8));
NOR2_X1 i_0_0_10 (.ZN (n_0_0_8), .A1 (n_0_0_6), .A2 (n_0_0_7));
INV_X1 i_0_0_9 (.ZN (n_0_0_7), .A (\i[2] ));
INV_X1 i_0_0_8 (.ZN (n_0_0_6), .A (\i[1] ));
OAI21_X1 i_0_0_7 (.ZN (n_0_0_5), .A (n_0_0_4), .B1 (\i[1] ), .B2 (\i[2] ));
INV_X1 i_0_0_6 (.ZN (n_0_0_4), .A (CLOCK_slh_n298));
NAND2_X1 i_0_0_5 (.ZN (n_0_0_3), .A1 (start_i[2]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_4 (.ZN (CLOCK_slh__n621), .A (n_0_0_2), .B1 (CLOCK_slh_n298), .B2 (\i[1] ));
NAND2_X1 i_0_0_3 (.ZN (n_0_0_2), .A1 (start_i[1]), .A2 (CLOCK_slh_n298));
OAI21_X1 i_0_0_2 (.ZN (CLOCK_slh__n623), .A (n_0_0_0), .B1 (n_0_0_1), .B2 (CLOCK_slh_n298));
INV_X1 i_0_0_1 (.ZN (n_0_0_1), .A (\i[0] ));
NAND2_X1 i_0_0_0 (.ZN (n_0_0_0), .A1 (start_i[0]), .A2 (CLOCK_slh_n298));
datapath__0_142 i_0_11 (.p_1 ({n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, n_0_229, 
    n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, n_0_223, n_0_222, n_0_221, n_0_220, 
    n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, 
    n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, 
    n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, 
    n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, 
    n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, 
    n_0_174, n_0_173, n_0_172, n_0_171}), .c ({\c[63] , \c[62] , \c[61] , \c[60] , 
    \c[59] , \c[58] , \c[57] , \c[56] , \c[55] , \c[54] , \c[53] , \c[52] , \c[51] , 
    \c[50] , \c[49] , \c[48] , \c[47] , \c[46] , \c[45] , \c[44] , \c[43] , \c[42] , 
    \c[41] , \c[40] , \c[39] , \c[38] , \c[37] , \c[36] , \c[35] , \c[34] , \c[33] , 
    \c[32] , \c[31] , \c[30] , \c[29] , \c[28] , \c[27] , \c[26] , \c[25] , \c[24] , 
    \c[23] , \c[22] , \c[21] , \c[20] , \c[19] , \c[18] , \c[17] , \c[16] , \c[15] , 
    \c[14] , \c[13] , \c[12] , \c[11] , \c[10] , \c[9] , \c[8] , \c[7] , \c[6] , 
    \c[5] , \c[4] , \c[3] , \c[2] , \c[1] , \c[0] }), .p_0 ({n_0_107, n_0_170, n_0_169, 
    n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, 
    n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, 
    n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, 
    n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, 
    n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, 
    n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, 
    n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108}));
datapath__0_128 i_0_4 (.p_0 ({uc_1, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
    n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, 
    n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
    n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, uc_2}), .p_1 ({1'b0 , \read_data2[31] , 
    \read_data2[30] , \read_data2[29] , \read_data2[28] , \read_data2[27] , \read_data2[26] , 
    \read_data2[25] , \read_data2[24] , \read_data2[23] , \read_data2[22] , \read_data2[21] , 
    \read_data2[20] , \read_data2[19] , \read_data2[18] , \read_data2[17] , \read_data2[16] , 
    \read_data2[15] , \read_data2[14] , \read_data2[13] , \read_data2[12] , \read_data2[11] , 
    \read_data2[10] , \read_data2[9] , \read_data2[8] , \read_data2[7] , \read_data2[6] , 
    \read_data2[5] , \read_data2[4] , \read_data2[3] , \read_data2[2] , \read_data2[1] , 
    \read_data2[0] }));
datapath i_0_3 (.p_0 ({n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, 
    n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
    n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, 
    n_0_6, n_0_5, n_0_4, uc_0}), .read_data2 ({\read_data2[31] , \read_data2[30] , 
    \read_data2[29] , \read_data2[28] , \read_data2[27] , \read_data2[26] , \read_data2[25] , 
    \read_data2[24] , \read_data2[23] , \read_data2[22] , \read_data2[21] , \read_data2[20] , 
    \read_data2[19] , \read_data2[18] , \read_data2[17] , \read_data2[16] , \read_data2[15] , 
    \read_data2[14] , \read_data2[13] , \read_data2[12] , \read_data2[11] , \read_data2[10] , 
    \read_data2[9] , \read_data2[8] , \read_data2[7] , \read_data2[6] , \read_data2[5] , 
    \read_data2[4] , \read_data2[3] , \read_data2[2] , \read_data2[1] , \read_data2[0] }));
DFF_X1 \res_reg[0]  (.Q (\res[0] ), .CK (CTS_n_tid0_68), .D (n_0_171));
DFF_X1 \res_reg[1]  (.Q (\res[1] ), .CK (CTS_n_tid0_68), .D (n_0_172));
DFF_X1 \res_reg[2]  (.Q (\res[2] ), .CK (CTS_n_tid0_68), .D (n_0_173));
DFF_X1 \res_reg[3]  (.Q (\res[3] ), .CK (CTS_n_tid0_68), .D (n_0_174));
DFF_X1 \res_reg[4]  (.Q (\res[4] ), .CK (CTS_n_tid0_68), .D (n_0_175));
DFF_X1 \res_reg[5]  (.Q (\res[5] ), .CK (CTS_n_tid0_68), .D (n_0_176));
DFF_X1 \res_reg[6]  (.Q (\res[6] ), .CK (CTS_n_tid0_68), .D (n_0_177));
DFF_X1 \res_reg[7]  (.Q (\res[7] ), .CK (CTS_n_tid0_68), .D (n_0_178));
DFF_X1 \res_reg[8]  (.Q (\res[8] ), .CK (CTS_n_tid0_68), .D (n_0_179));
DFF_X1 \res_reg[9]  (.Q (\res[9] ), .CK (CTS_n_tid0_68), .D (n_0_180));
DFF_X1 \res_reg[10]  (.Q (\res[10] ), .CK (CTS_n_tid0_68), .D (n_0_181));
DFF_X1 \res_reg[11]  (.Q (\res[11] ), .CK (CTS_n_tid0_68), .D (n_0_182));
DFF_X1 \res_reg[12]  (.Q (\res[12] ), .CK (CTS_n_tid0_68), .D (n_0_183));
DFF_X1 \res_reg[13]  (.Q (\res[13] ), .CK (CTS_n_tid0_68), .D (n_0_184));
DFF_X1 \res_reg[14]  (.Q (\res[14] ), .CK (CTS_n_tid0_68), .D (n_0_185));
DFF_X1 \res_reg[15]  (.Q (\res[15] ), .CK (CTS_n_tid0_68), .D (n_0_186));
DFF_X1 \res_reg[16]  (.Q (\res[16] ), .CK (CTS_n_tid0_68), .D (n_0_187));
DFF_X1 \res_reg[17]  (.Q (\res[17] ), .CK (CTS_n_tid0_68), .D (n_0_188));
DFF_X1 \res_reg[18]  (.Q (\res[18] ), .CK (CTS_n_tid0_68), .D (n_0_189));
DFF_X1 \res_reg[19]  (.Q (\res[19] ), .CK (CTS_n_tid0_68), .D (n_0_190));
DFF_X1 \res_reg[20]  (.Q (\res[20] ), .CK (CTS_n_tid0_68), .D (n_0_191));
DFF_X1 \res_reg[21]  (.Q (\res[21] ), .CK (CTS_n_tid0_68), .D (n_0_192));
DFF_X1 \res_reg[22]  (.Q (\res[22] ), .CK (CTS_n_tid0_68), .D (n_0_193));
DFF_X1 \res_reg[23]  (.Q (\res[23] ), .CK (CTS_n_tid0_68), .D (n_0_194));
DFF_X1 \res_reg[24]  (.Q (\res[24] ), .CK (CTS_n_tid0_68), .D (n_0_195));
DFF_X1 \res_reg[25]  (.Q (\res[25] ), .CK (CTS_n_tid0_68), .D (n_0_196));
DFF_X1 \res_reg[26]  (.Q (\res[26] ), .CK (CTS_n_tid0_68), .D (n_0_197));
DFF_X1 \res_reg[27]  (.Q (\res[27] ), .CK (CTS_n_tid0_68), .D (n_0_198));
DFF_X1 \res_reg[28]  (.Q (\res[28] ), .CK (CTS_n_tid0_68), .D (n_0_199));
DFF_X1 \res_reg[29]  (.Q (\res[29] ), .CK (CTS_n_tid0_68), .D (n_0_200));
DFF_X1 \res_reg[30]  (.Q (\res[30] ), .CK (CTS_n_tid0_68), .D (n_0_201));
DFF_X1 \res_reg[31]  (.Q (\res[31] ), .CK (CTS_n_tid0_68), .D (n_0_202));
DFF_X1 \res_reg[32]  (.Q (\res[32] ), .CK (CTS_n_tid0_68), .D (n_0_203));
DFF_X1 \res_reg[33]  (.Q (\res[33] ), .CK (CTS_n_tid0_68), .D (n_0_204));
DFF_X1 \res_reg[34]  (.Q (\res[34] ), .CK (CTS_n_tid0_68), .D (n_0_205));
DFF_X1 \res_reg[35]  (.Q (\res[35] ), .CK (CTS_n_tid0_68), .D (n_0_206));
DFF_X1 \res_reg[36]  (.Q (\res[36] ), .CK (CTS_n_tid0_68), .D (n_0_207));
DFF_X1 \res_reg[37]  (.Q (\res[37] ), .CK (CTS_n_tid0_68), .D (n_0_208));
DFF_X1 \res_reg[38]  (.Q (\res[38] ), .CK (CTS_n_tid0_68), .D (n_0_209));
DFF_X1 \res_reg[39]  (.Q (\res[39] ), .CK (CTS_n_tid0_68), .D (n_0_210));
DFF_X1 \res_reg[40]  (.Q (\res[40] ), .CK (CTS_n_tid0_68), .D (n_0_211));
DFF_X1 \res_reg[41]  (.Q (\res[41] ), .CK (CTS_n_tid0_68), .D (n_0_212));
DFF_X1 \res_reg[42]  (.Q (\res[42] ), .CK (CTS_n_tid0_68), .D (n_0_213));
DFF_X1 \res_reg[43]  (.Q (\res[43] ), .CK (CTS_n_tid0_68), .D (n_0_214));
DFF_X1 \res_reg[44]  (.Q (\res[44] ), .CK (CTS_n_tid0_68), .D (n_0_215));
DFF_X1 \res_reg[45]  (.Q (\res[45] ), .CK (CTS_n_tid0_68), .D (n_0_216));
DFF_X1 \res_reg[46]  (.Q (\res[46] ), .CK (CTS_n_tid0_68), .D (n_0_217));
DFF_X1 \res_reg[47]  (.Q (\res[47] ), .CK (CTS_n_tid0_68), .D (n_0_218));
DFF_X1 \res_reg[48]  (.Q (\res[48] ), .CK (CTS_n_tid0_68), .D (n_0_219));
DFF_X1 \res_reg[49]  (.Q (\res[49] ), .CK (CTS_n_tid0_68), .D (n_0_220));
DFF_X1 \res_reg[50]  (.Q (\res[50] ), .CK (CTS_n_tid0_68), .D (n_0_221));
DFF_X1 \res_reg[51]  (.Q (\res[51] ), .CK (CTS_n_tid0_68), .D (n_0_222));
DFF_X1 \res_reg[52]  (.Q (\res[52] ), .CK (CTS_n_tid0_68), .D (n_0_223));
DFF_X1 \res_reg[53]  (.Q (\res[53] ), .CK (CTS_n_tid0_68), .D (n_0_224));
DFF_X1 \res_reg[54]  (.Q (\res[54] ), .CK (CTS_n_tid0_68), .D (n_0_225));
DFF_X1 \res_reg[55]  (.Q (\res[55] ), .CK (CTS_n_tid0_68), .D (n_0_226));
DFF_X1 \res_reg[56]  (.Q (\res[56] ), .CK (CTS_n_tid0_68), .D (n_0_227));
DFF_X1 \res_reg[57]  (.Q (\res[57] ), .CK (CTS_n_tid0_68), .D (n_0_228));
DFF_X1 \res_reg[58]  (.Q (\res[58] ), .CK (CTS_n_tid0_68), .D (n_0_229));
DFF_X1 \res_reg[59]  (.Q (\res[59] ), .CK (CTS_n_tid0_68), .D (n_0_230));
DFF_X1 \res_reg[60]  (.Q (\res[60] ), .CK (CTS_n_tid0_68), .D (n_0_231));
DFF_X1 \res_reg[61]  (.Q (\res[61] ), .CK (CTS_n_tid0_68), .D (n_0_232));
DFF_X1 \res_reg[62]  (.Q (\res[62] ), .CK (CTS_n_tid0_68), .D (n_0_233));
DFF_X1 \res_reg[63]  (.Q (\res[63] ), .CK (CTS_n_tid0_68), .D (n_0_234));
CLKGATETST_X8 clk_gate_res_reg (.GCK (CTS_n_tid0_69), .CK (CTS_n_tid1_199), .E (hfn_ipo_n41), .SE (1'b0 ));
regFile64 r2 (.read_data ({read_data3[63], read_data3[62], read_data3[61], read_data3[60], 
    read_data3[59], read_data3[58], read_data3[57], read_data3[56], read_data3[55], 
    read_data3[54], read_data3[53], read_data3[52], read_data3[51], read_data3[50], 
    read_data3[49], read_data3[48], read_data3[47], read_data3[46], read_data3[45], 
    read_data3[44], read_data3[43], read_data3[42], read_data3[41], read_data3[40], 
    read_data3[39], read_data3[38], read_data3[37], read_data3[36], read_data3[35], 
    read_data3[34], read_data3[33], read_data3[32], read_data3[31], read_data3[30], 
    read_data3[29], read_data3[28], read_data3[27], read_data3[26], read_data3[25], 
    read_data3[24], read_data3[23], read_data3[22], read_data3[21], read_data3[20], 
    read_data3[19], read_data3[18], read_data3[17], read_data3[16], read_data3[15], 
    read_data3[14], read_data3[13], read_data3[12], read_data3[11], read_data3[10], 
    read_data3[9], read_data3[8], read_data3[7], read_data3[6], read_data3[5], read_data3[4], 
    read_data3[3], read_data3[2], read_data3[1], read_data3[0]}), .write_data ({\res[63] , 
    \res[62] , \res[61] , \res[60] , \res[59] , \res[58] , \res[57] , \res[56] , 
    \res[55] , \res[54] , \res[53] , \res[52] , \res[51] , \res[50] , \res[49] , 
    \res[48] , \res[47] , \res[46] , \res[45] , \res[44] , \res[43] , \res[42] , 
    \res[41] , \res[40] , \res[39] , \res[38] , \res[37] , \res[36] , \res[35] , 
    \res[34] , \res[33] , \res[32] , \res[31] , \res[30] , \res[29] , \res[28] , 
    \res[27] , \res[26] , \res[25] , \res[24] , \res[23] , \res[22] , \res[21] , 
    \res[20] , \res[19] , \res[18] , \res[17] , \res[16] , \res[15] , \res[14] , 
    \res[13] , \res[12] , \res[11] , \res[10] , \res[9] , \res[8] , \res[7] , \res[6] , 
    \res[5] , \res[4] , \res[3] , \res[2] , \res[1] , \res[0] }), .clk__CTS_1_PP_0 (CTS_n_tid1_188));
regFile r (.read_data2 ({\read_data2[31] , \read_data2[30] , \read_data2[29] , \read_data2[28] , 
    \read_data2[27] , \read_data2[26] , \read_data2[25] , \read_data2[24] , \read_data2[23] , 
    \read_data2[22] , \read_data2[21] , \read_data2[20] , \read_data2[19] , \read_data2[18] , 
    \read_data2[17] , \read_data2[16] , \read_data2[15] , \read_data2[14] , \read_data2[13] , 
    \read_data2[12] , \read_data2[11] , \read_data2[10] , \read_data2[9] , \read_data2[8] , 
    \read_data2[7] , \read_data2[6] , \read_data2[5] , \read_data2[4] , \read_data2[3] , 
    \read_data2[2] , \read_data2[1] , \read_data2[0] }), .read_data ({\read_data[31] , 
    \read_data[30] , \read_data[29] , \read_data[28] , \read_data[27] , \read_data[26] , 
    \read_data[25] , \read_data[24] , \read_data[23] , \read_data[22] , \read_data[21] , 
    \read_data[20] , \read_data[19] , \read_data[18] , \read_data[17] , \read_data[16] , 
    \read_data[15] , \read_data[14] , \read_data[13] , \read_data[12] , \read_data[11] , 
    \read_data[10] , \read_data[9] , \read_data[8] , \read_data[7] , \read_data[6] , 
    \read_data[5] , \read_data[4] , \read_data[3] , \read_data[2] , \read_data[1] , 
    \read_data[0] }), .clk__CTS_1_PP_0 (CTS_n_tid1_188), .clk__CTS_1_PP_3 (CTS_n_tid1_199)
    , .write_data2 ({CLOCK_slh_n363, CLOCK_slh_n558, CLOCK_slh_n553, CLOCK_slh_n548, 
    CLOCK_slh_n358, CLOCK_slh_n543, CLOCK_slh_n538, CLOCK_slh_n533, CLOCK_slh_n528, 
    CLOCK_slh_n408, CLOCK_slh_n523, CLOCK_slh_n518, CLOCK_slh_n513, CLOCK_slh_n403, 
    CLOCK_slh_n573, CLOCK_slh_n618, CLOCK_slh_n508, CLOCK_slh_n373, CLOCK_slh_n503, 
    CLOCK_slh_n498, CLOCK_slh_n398, CLOCK_slh_n493, CLOCK_slh_n568, CLOCK_slh_n413, 
    CLOCK_slh_n563, CLOCK_slh_n378, CLOCK_slh_n608, CLOCK_slh_n598, CLOCK_slh_n333, 
    CLOCK_slh_n303, CLOCK_slh_n323, CLOCK_slh_n318}), .write_data ({CLOCK_slh_n313, 
    CLOCK_slh_n338, CLOCK_slh_n478, CLOCK_slh_n383, CLOCK_slh_n473, CLOCK_slh_n468, 
    CLOCK_slh_n463, CLOCK_slh_n353, CLOCK_slh_n458, CLOCK_slh_n453, CLOCK_slh_n588, 
    CLOCK_slh_n448, CLOCK_slh_n438, CLOCK_slh_n583, CLOCK_slh_n433, CLOCK_slh_n348, 
    CLOCK_slh_n308, CLOCK_slh_n428, CLOCK_slh_n613, CLOCK_slh_n423, CLOCK_slh_n343, 
    CLOCK_slh_n578, CLOCK_slh_n368, CLOCK_slh_n603, CLOCK_slh_n418, CLOCK_slh_n488, 
    CLOCK_slh_n393, CLOCK_slh_n388, CLOCK_slh_n483, CLOCK_slh_n593, CLOCK_slh_n443, 
    CLOCK_slh_n328}), .write_en (write_en), .clk__CTS_1_PP_4 (clk));
CLKBUF_X2 hfn_ipo_c49 (.Z (hfn_ipo_n49), .A (\shift[0] ));
CLKBUF_X2 hfn_ipo_c50 (.Z (hfn_ipo_n50), .A (\shift[0] ));
BUF_X4 hfn_ipo_c41 (.Z (hfn_ipo_n41), .A (n_0_105));
CLKBUF_X3 CTS_L3_c_tid0_69 (.Z (CTS_n_tid0_68), .A (CTS_n_tid0_69));
CLKBUF_X2 hfn_ipo_c45 (.Z (hfn_ipo_n45), .A (\shift[2] ));
CLKBUF_X1 hfn_ipo_c46 (.Z (hfn_ipo_n46), .A (\shift[2] ));
CLKBUF_X2 hfn_ipo_c35 (.Z (hfn_ipo_n35), .A (n_0_0_19));
CLKBUF_X1 hfn_ipo_c36 (.Z (hfn_ipo_n36), .A (n_0_0_19));
CLKBUF_X1 hfn_ipo_c37 (.Z (hfn_ipo_n37), .A (n_0_0_23));
CLKBUF_X2 CTS_L3_c_tid1_133 (.Z (CTS_n_tid1_147), .A (CTS_n_tid1_188));
CLKBUF_X1 CLOCK_slh__c209 (.Z (CLOCK_slh_n298), .A (start));
BUF_X4 hfn_ipo_c43 (.Z (hfn_ipo_n43), .A (n_0_0_38));
CLKBUF_X1 hfn_ipo_c44 (.Z (hfn_ipo_n44), .A (n_0_0_38));
CLKBUF_X1 hfn_ipo_c47 (.Z (hfn_ipo_n47), .A (\shift[1] ));
CLKBUF_X1 hfn_ipo_c48 (.Z (hfn_ipo_n48), .A (\shift[1] ));
BUF_X4 drc_ipo_c51 (.Z (drc_ipo_n51), .A (n_0_0_192));
CLKBUF_X2 hfn_ipo_c39 (.Z (hfn_ipo_n39), .A (n_0_0_24));
CLKBUF_X1 CLOCK_slh__c211 (.Z (CLOCK_slh__n699), .A (b[2]));
CLKBUF_X1 CLOCK_slh__c215 (.Z (CLOCK_slh__n999), .A (a[31]));
CLKBUF_X1 CLOCK_slh__c213 (.Z (CLOCK_slh__n921), .A (a[15]));
CLKBUF_X1 CLOCK_slh__c217 (.Z (CLOCK_slh__n639), .A (b[0]));
CLKBUF_X1 CLOCK_slh__c225 (.Z (CLOCK_slh__n819), .A (a[30]));
CLKBUF_X1 CLOCK_slh__c227 (.Z (CLOCK_slh__n717), .A (a[11]));
CLKBUF_X1 CLOCK_slh__c219 (.Z (CLOCK_slh__n975), .A (b[1]));
CLKBUF_X1 CLOCK_slh__c221 (.Z (CLOCK_slh__n807), .A (a[0]));
CLKBUF_X1 CLOCK_slh__c223 (.Z (CLOCK_slh__n801), .A (b[3]));
CLKBUF_X2 CTS_L3_c_tid1_189 (.Z (CTS_n_tid1_187), .A (CTS_n_tid1_188));
CLKBUF_X1 CLOCK_slh__c229 (.Z (CLOCK_slh__n711), .A (a[16]));
CLKBUF_X1 CLOCK_slh__c231 (.Z (CLOCK_slh__n705), .A (a[24]));
CLKBUF_X1 CLOCK_slh__c233 (.Z (CLOCK_slh__n723), .A (b[27]));
CLKBUF_X1 CLOCK_slh__c235 (.Z (CLOCK_slh__n729), .A (b[31]));
CLKBUF_X1 CLOCK_slh__c237 (.Z (CLOCK_slh__n1011), .A (a[9]));
CLKBUF_X1 CLOCK_slh__c239 (.Z (CLOCK_slh__n765), .A (b[14]));
CLKBUF_X1 CLOCK_slh__c241 (.Z (CLOCK_slh__n771), .A (b[6]));
CLKBUF_X1 CLOCK_slh__c243 (.Z (CLOCK_slh__n777), .A (a[28]));
CLKBUF_X1 CLOCK_slh__c245 (.Z (CLOCK_slh__n783), .A (a[4]));
CLKBUF_X1 CLOCK_slh__c247 (.Z (CLOCK_slh__n759), .A (a[5]));
CLKBUF_X1 CLOCK_slh__c249 (.Z (CLOCK_slh__n645), .A (b[11]));
CLKBUF_X1 CLOCK_slh__c251 (.Z (CLOCK_slh__n735), .A (b[18]));
CLKBUF_X1 CLOCK_slh__c253 (.Z (CLOCK_slh__n651), .A (b[22]));
CLKBUF_X1 CLOCK_slh__c255 (.Z (CLOCK_slh__n789), .A (b[8]));
CLKBUF_X1 CLOCK_slh__c257 (.Z (CLOCK_slh__n795), .A (a[7]));
CLKBUF_X1 CLOCK_slh__c259 (.Z (CLOCK_slh__n741), .A (a[12]));
CLKBUF_X1 CLOCK_slh__c261 (.Z (CLOCK_slh__n993), .A (a[14]));
CLKBUF_X1 CLOCK_slh__c263 (.Z (CLOCK_slh__n1017), .A (a[17]));
CLKBUF_X1 CLOCK_slh__c265 (.Z (CLOCK_slh__n825), .A (a[19]));
CLKBUF_X1 CLOCK_slh__c267 (.Z (CLOCK_slh__n981), .A (a[1]));
CLKBUF_X1 CLOCK_slh__c269 (.Z (CLOCK_slh__n753), .A (a[20]));
CLKBUF_X1 CLOCK_slh__c271 (.Z (CLOCK_slh__n969), .A (a[22]));
CLKBUF_X1 CLOCK_slh__c273 (.Z (CLOCK_slh__n903), .A (a[23]));
CLKBUF_X1 CLOCK_slh__c275 (.Z (CLOCK_slh__n657), .A (a[25]));
CLKBUF_X1 CLOCK_slh__c277 (.Z (CLOCK_slh__n873), .A (a[26]));
CLKBUF_X1 CLOCK_slh__c279 (.Z (CLOCK_slh__n681), .A (a[27]));
CLKBUF_X1 CLOCK_slh__c281 (.Z (CLOCK_slh__n867), .A (a[29]));
CLKBUF_X1 CLOCK_slh__c283 (.Z (CLOCK_slh__n693), .A (a[3]));
CLKBUF_X1 CLOCK_slh__c285 (.Z (CLOCK_slh__n927), .A (a[6]));
CLKBUF_X1 CLOCK_slh__c287 (.Z (CLOCK_slh__n891), .A (b[10]));
CLKBUF_X1 CLOCK_slh__c289 (.Z (CLOCK_slh__n669), .A (b[12]));
CLKBUF_X1 CLOCK_slh__c291 (.Z (CLOCK_slh__n909), .A (b[13]));
CLKBUF_X1 CLOCK_slh__c293 (.Z (CLOCK_slh__n675), .A (b[15]));
CLKBUF_X1 CLOCK_slh__c295 (.Z (CLOCK_slh__n879), .A (b[19]));
CLKBUF_X1 CLOCK_slh__c297 (.Z (CLOCK_slh__n687), .A (b[20]));
CLKBUF_X1 CLOCK_slh__c299 (.Z (CLOCK_slh__n897), .A (b[21]));
CLKBUF_X1 CLOCK_slh__c301 (.Z (CLOCK_slh__n837), .A (b[23]));
CLKBUF_X1 CLOCK_slh__c303 (.Z (CLOCK_slh__n933), .A (b[24]));
CLKBUF_X1 CLOCK_slh__c305 (.Z (CLOCK_slh__n747), .A (b[25]));
CLKBUF_X1 CLOCK_slh__c307 (.Z (CLOCK_slh__n1005), .A (b[26]));
CLKBUF_X1 CLOCK_slh__c309 (.Z (CLOCK_slh__n663), .A (b[28]));
CLKBUF_X1 CLOCK_slh__c311 (.Z (CLOCK_slh__n963), .A (b[29]));
CLKBUF_X1 CLOCK_slh__c313 (.Z (CLOCK_slh__n831), .A (b[30]));
CLKBUF_X1 CLOCK_slh__c315 (.Z (CLOCK_slh__n813), .A (b[7]));
CLKBUF_X1 CLOCK_slh__c317 (.Z (CLOCK_slh__n843), .A (b[9]));
CLKBUF_X1 CLOCK_slh__c319 (.Z (CLOCK_slh__n915), .A (b[17]));
CLKBUF_X1 CLOCK_slh__c321 (.Z (CLOCK_slh__n855), .A (a[10]));
CLKBUF_X1 CLOCK_slh__c323 (.Z (CLOCK_slh__n861), .A (a[18]));
CLKBUF_X1 CLOCK_slh__c325 (.Z (CLOCK_slh__n885), .A (a[21]));
CLKBUF_X1 CLOCK_slh__c327 (.Z (CLOCK_slh__n849), .A (a[2]));
CLKBUF_X1 CLOCK_slh__c329 (.Z (CLOCK_slh__n939), .A (b[4]));
CLKBUF_X1 CLOCK_slh__c331 (.Z (CLOCK_slh__n945), .A (a[8]));
CLKBUF_X1 CLOCK_slh__c333 (.Z (CLOCK_slh__n951), .A (b[5]));
CLKBUF_X1 CLOCK_slh__c335 (.Z (CLOCK_slh__n987), .A (a[13]));
CLKBUF_X1 CLOCK_slh__c337 (.Z (CLOCK_slh__n957), .A (b[16]));
CLKBUF_X1 CLOCK_slh__c339 (.Z (n_0_71), .A (CLOCK_slh__n619));
CLKBUF_X1 CLOCK_slh__c341 (.Z (n_0_2), .A (CLOCK_slh__n621));
CLKBUF_X1 CLOCK_slh__c343 (.Z (n_0_1), .A (CLOCK_slh__n623));
CLKBUF_X1 CLOCK_slh__c345 (.Z (n_0_70), .A (CLOCK_slh__n625));
CLKBUF_X1 CLOCK_slh__c347 (.Z (n_0_66), .A (CLOCK_slh__n627));
CLKBUF_X1 CLOCK_slh__c349 (.Z (n_0_3), .A (CLOCK_slh__n629));
CLKBUF_X1 CLOCK_slh__c351 (.Z (n_0_67), .A (CLOCK_slh__n631));
CLKBUF_X1 CLOCK_slh__c353 (.Z (n_0_73), .A (CLOCK_slh__n633));
CLKBUF_X1 CLOCK_slh__c355 (.Z (n_0_74), .A (CLOCK_slh__n635));
CLKBUF_X1 CLOCK_slh__c357 (.Z (n_0_72), .A (CLOCK_slh__n637));
CLKBUF_X1 CLOCK_slh__c359 (.Z (CLOCK_slh__n640), .A (CLOCK_slh__n639));
CLKBUF_X1 CLOCK_slh__c360 (.Z (CLOCK_slh__n641), .A (CLOCK_slh__n640));
CLKBUF_X1 CLOCK_slh__c361 (.Z (CLOCK_slh_n318), .A (CLOCK_slh__n641));
CLKBUF_X1 CLOCK_slh__c365 (.Z (CLOCK_slh__n646), .A (CLOCK_slh__n645));
CLKBUF_X1 CLOCK_slh__c366 (.Z (CLOCK_slh__n647), .A (CLOCK_slh__n646));
CLKBUF_X1 CLOCK_slh__c367 (.Z (CLOCK_slh_n398), .A (CLOCK_slh__n647));
CLKBUF_X1 CLOCK_slh__c371 (.Z (CLOCK_slh__n652), .A (CLOCK_slh__n651));
CLKBUF_X1 CLOCK_slh__c372 (.Z (CLOCK_slh__n653), .A (CLOCK_slh__n652));
CLKBUF_X1 CLOCK_slh__c373 (.Z (CLOCK_slh_n408), .A (CLOCK_slh__n653));
CLKBUF_X1 CLOCK_slh__c377 (.Z (CLOCK_slh__n658), .A (CLOCK_slh__n657));
CLKBUF_X1 CLOCK_slh__c378 (.Z (CLOCK_slh__n659), .A (CLOCK_slh__n658));
CLKBUF_X1 CLOCK_slh__c379 (.Z (CLOCK_slh_n463), .A (CLOCK_slh__n659));
CLKBUF_X1 CLOCK_slh__c383 (.Z (CLOCK_slh__n664), .A (CLOCK_slh__n663));
CLKBUF_X1 CLOCK_slh__c384 (.Z (CLOCK_slh__n665), .A (CLOCK_slh__n664));
CLKBUF_X1 CLOCK_slh__c385 (.Z (CLOCK_slh_n548), .A (CLOCK_slh__n665));
CLKBUF_X1 CLOCK_slh__c389 (.Z (CLOCK_slh__n670), .A (CLOCK_slh__n669));
CLKBUF_X1 CLOCK_slh__c390 (.Z (CLOCK_slh__n671), .A (CLOCK_slh__n670));
CLKBUF_X1 CLOCK_slh__c391 (.Z (CLOCK_slh_n498), .A (CLOCK_slh__n671));
CLKBUF_X1 CLOCK_slh__c395 (.Z (CLOCK_slh__n676), .A (CLOCK_slh__n675));
CLKBUF_X1 CLOCK_slh__c396 (.Z (CLOCK_slh__n677), .A (CLOCK_slh__n676));
CLKBUF_X1 CLOCK_slh__c397 (.Z (CLOCK_slh_n508), .A (CLOCK_slh__n677));
CLKBUF_X1 CLOCK_slh__c401 (.Z (CLOCK_slh__n682), .A (CLOCK_slh__n681));
CLKBUF_X1 CLOCK_slh__c402 (.Z (CLOCK_slh__n683), .A (CLOCK_slh__n682));
CLKBUF_X1 CLOCK_slh__c403 (.Z (CLOCK_slh_n473), .A (CLOCK_slh__n683));
CLKBUF_X1 CLOCK_slh__c407 (.Z (CLOCK_slh__n688), .A (CLOCK_slh__n687));
CLKBUF_X1 CLOCK_slh__c408 (.Z (CLOCK_slh__n689), .A (CLOCK_slh__n688));
CLKBUF_X1 CLOCK_slh__c409 (.Z (CLOCK_slh_n518), .A (CLOCK_slh__n689));
CLKBUF_X1 CLOCK_slh__c413 (.Z (CLOCK_slh__n694), .A (CLOCK_slh__n693));
CLKBUF_X1 CLOCK_slh__c414 (.Z (CLOCK_slh__n695), .A (CLOCK_slh__n694));
CLKBUF_X1 CLOCK_slh__c415 (.Z (CLOCK_slh_n483), .A (CLOCK_slh__n695));
CLKBUF_X1 CLOCK_slh__c419 (.Z (CLOCK_slh__n700), .A (CLOCK_slh__n699));
CLKBUF_X1 CLOCK_slh__c420 (.Z (CLOCK_slh__n701), .A (CLOCK_slh__n700));
CLKBUF_X1 CLOCK_slh__c421 (.Z (CLOCK_slh_n303), .A (CLOCK_slh__n701));
CLKBUF_X1 CLOCK_slh__c425 (.Z (CLOCK_slh__n706), .A (CLOCK_slh__n705));
CLKBUF_X1 CLOCK_slh__c426 (.Z (CLOCK_slh__n707), .A (CLOCK_slh__n706));
CLKBUF_X1 CLOCK_slh__c427 (.Z (CLOCK_slh_n353), .A (CLOCK_slh__n707));
CLKBUF_X1 CLOCK_slh__c431 (.Z (CLOCK_slh__n712), .A (CLOCK_slh__n711));
CLKBUF_X1 CLOCK_slh__c432 (.Z (CLOCK_slh__n713), .A (CLOCK_slh__n712));
CLKBUF_X1 CLOCK_slh__c433 (.Z (CLOCK_slh_n348), .A (CLOCK_slh__n713));
CLKBUF_X1 CLOCK_slh__c437 (.Z (CLOCK_slh__n718), .A (CLOCK_slh__n717));
CLKBUF_X1 CLOCK_slh__c438 (.Z (CLOCK_slh__n719), .A (CLOCK_slh__n718));
CLKBUF_X1 CLOCK_slh__c439 (.Z (CLOCK_slh_n343), .A (CLOCK_slh__n719));
CLKBUF_X1 CLOCK_slh__c443 (.Z (CLOCK_slh__n724), .A (CLOCK_slh__n723));
CLKBUF_X1 CLOCK_slh__c444 (.Z (CLOCK_slh__n725), .A (CLOCK_slh__n724));
CLKBUF_X1 CLOCK_slh__c445 (.Z (CLOCK_slh_n358), .A (CLOCK_slh__n725));
CLKBUF_X1 CLOCK_slh__c449 (.Z (CLOCK_slh__n730), .A (CLOCK_slh__n729));
CLKBUF_X1 CLOCK_slh__c450 (.Z (CLOCK_slh__n731), .A (CLOCK_slh__n730));
CLKBUF_X1 CLOCK_slh__c451 (.Z (CLOCK_slh_n363), .A (CLOCK_slh__n731));
CLKBUF_X1 CLOCK_slh__c455 (.Z (CLOCK_slh__n736), .A (CLOCK_slh__n735));
CLKBUF_X1 CLOCK_slh__c456 (.Z (CLOCK_slh__n737), .A (CLOCK_slh__n736));
CLKBUF_X1 CLOCK_slh__c457 (.Z (CLOCK_slh_n403), .A (CLOCK_slh__n737));
CLKBUF_X1 CLOCK_slh__c461 (.Z (CLOCK_slh__n742), .A (CLOCK_slh__n741));
CLKBUF_X1 CLOCK_slh__c462 (.Z (CLOCK_slh__n743), .A (CLOCK_slh__n742));
CLKBUF_X1 CLOCK_slh__c463 (.Z (CLOCK_slh_n423), .A (CLOCK_slh__n743));
CLKBUF_X1 CLOCK_slh__c467 (.Z (CLOCK_slh__n748), .A (CLOCK_slh__n747));
CLKBUF_X1 CLOCK_slh__c468 (.Z (CLOCK_slh__n749), .A (CLOCK_slh__n748));
CLKBUF_X1 CLOCK_slh__c469 (.Z (CLOCK_slh_n538), .A (CLOCK_slh__n749));
CLKBUF_X1 CLOCK_slh__c473 (.Z (CLOCK_slh__n754), .A (CLOCK_slh__n753));
CLKBUF_X1 CLOCK_slh__c474 (.Z (CLOCK_slh__n755), .A (CLOCK_slh__n754));
CLKBUF_X1 CLOCK_slh__c475 (.Z (CLOCK_slh_n448), .A (CLOCK_slh__n755));
CLKBUF_X1 CLOCK_slh__c479 (.Z (CLOCK_slh__n760), .A (CLOCK_slh__n759));
CLKBUF_X1 CLOCK_slh__c480 (.Z (CLOCK_slh__n761), .A (CLOCK_slh__n760));
CLKBUF_X1 CLOCK_slh__c481 (.Z (CLOCK_slh_n393), .A (CLOCK_slh__n761));
CLKBUF_X1 CLOCK_slh__c485 (.Z (CLOCK_slh__n766), .A (CLOCK_slh__n765));
CLKBUF_X1 CLOCK_slh__c486 (.Z (CLOCK_slh__n767), .A (CLOCK_slh__n766));
CLKBUF_X1 CLOCK_slh__c487 (.Z (CLOCK_slh_n373), .A (CLOCK_slh__n767));
CLKBUF_X1 CLOCK_slh__c491 (.Z (CLOCK_slh__n772), .A (CLOCK_slh__n771));
CLKBUF_X1 CLOCK_slh__c492 (.Z (CLOCK_slh__n773), .A (CLOCK_slh__n772));
CLKBUF_X1 CLOCK_slh__c493 (.Z (CLOCK_slh_n378), .A (CLOCK_slh__n773));
CLKBUF_X1 CLOCK_slh__c497 (.Z (CLOCK_slh__n778), .A (CLOCK_slh__n777));
CLKBUF_X1 CLOCK_slh__c498 (.Z (CLOCK_slh__n779), .A (CLOCK_slh__n778));
CLKBUF_X1 CLOCK_slh__c499 (.Z (CLOCK_slh_n383), .A (CLOCK_slh__n779));
CLKBUF_X1 CLOCK_slh__c503 (.Z (CLOCK_slh__n784), .A (CLOCK_slh__n783));
CLKBUF_X1 CLOCK_slh__c504 (.Z (CLOCK_slh__n785), .A (CLOCK_slh__n784));
CLKBUF_X1 CLOCK_slh__c505 (.Z (CLOCK_slh_n388), .A (CLOCK_slh__n785));
CLKBUF_X1 CLOCK_slh__c509 (.Z (CLOCK_slh__n790), .A (CLOCK_slh__n789));
CLKBUF_X1 CLOCK_slh__c510 (.Z (CLOCK_slh__n791), .A (CLOCK_slh__n790));
CLKBUF_X1 CLOCK_slh__c511 (.Z (CLOCK_slh_n413), .A (CLOCK_slh__n791));
CLKBUF_X1 CLOCK_slh__c515 (.Z (CLOCK_slh__n796), .A (CLOCK_slh__n795));
CLKBUF_X1 CLOCK_slh__c516 (.Z (CLOCK_slh__n797), .A (CLOCK_slh__n796));
CLKBUF_X1 CLOCK_slh__c517 (.Z (CLOCK_slh_n418), .A (CLOCK_slh__n797));
CLKBUF_X1 CLOCK_slh__c521 (.Z (CLOCK_slh__n802), .A (CLOCK_slh__n801));
CLKBUF_X1 CLOCK_slh__c522 (.Z (CLOCK_slh__n803), .A (CLOCK_slh__n802));
CLKBUF_X1 CLOCK_slh__c523 (.Z (CLOCK_slh_n333), .A (CLOCK_slh__n803));
CLKBUF_X1 CLOCK_slh__c527 (.Z (CLOCK_slh__n808), .A (CLOCK_slh__n807));
CLKBUF_X1 CLOCK_slh__c528 (.Z (CLOCK_slh__n809), .A (CLOCK_slh__n808));
CLKBUF_X1 CLOCK_slh__c529 (.Z (CLOCK_slh_n328), .A (CLOCK_slh__n809));
CLKBUF_X1 CLOCK_slh__c533 (.Z (CLOCK_slh__n814), .A (CLOCK_slh__n813));
CLKBUF_X1 CLOCK_slh__c534 (.Z (CLOCK_slh__n815), .A (CLOCK_slh__n814));
CLKBUF_X1 CLOCK_slh__c535 (.Z (CLOCK_slh_n563), .A (CLOCK_slh__n815));
CLKBUF_X1 CLOCK_slh__c539 (.Z (CLOCK_slh__n820), .A (CLOCK_slh__n819));
CLKBUF_X1 CLOCK_slh__c540 (.Z (CLOCK_slh__n821), .A (CLOCK_slh__n820));
CLKBUF_X1 CLOCK_slh__c541 (.Z (CLOCK_slh_n338), .A (CLOCK_slh__n821));
CLKBUF_X1 CLOCK_slh__c545 (.Z (CLOCK_slh__n826), .A (CLOCK_slh__n825));
CLKBUF_X1 CLOCK_slh__c546 (.Z (CLOCK_slh__n827), .A (CLOCK_slh__n826));
CLKBUF_X1 CLOCK_slh__c547 (.Z (CLOCK_slh_n438), .A (CLOCK_slh__n827));
CLKBUF_X1 CLOCK_slh__c551 (.Z (CLOCK_slh__n832), .A (CLOCK_slh__n831));
CLKBUF_X1 CLOCK_slh__c552 (.Z (CLOCK_slh__n833), .A (CLOCK_slh__n832));
CLKBUF_X1 CLOCK_slh__c553 (.Z (CLOCK_slh_n558), .A (CLOCK_slh__n833));
CLKBUF_X1 CLOCK_slh__c557 (.Z (CLOCK_slh__n838), .A (CLOCK_slh__n837));
CLKBUF_X1 CLOCK_slh__c558 (.Z (CLOCK_slh__n839), .A (CLOCK_slh__n838));
CLKBUF_X1 CLOCK_slh__c559 (.Z (CLOCK_slh_n528), .A (CLOCK_slh__n839));
CLKBUF_X1 CLOCK_slh__c563 (.Z (CLOCK_slh__n844), .A (CLOCK_slh__n843));
CLKBUF_X1 CLOCK_slh__c564 (.Z (CLOCK_slh__n845), .A (CLOCK_slh__n844));
CLKBUF_X1 CLOCK_slh__c565 (.Z (CLOCK_slh_n568), .A (CLOCK_slh__n845));
CLKBUF_X1 CLOCK_slh__c569 (.Z (CLOCK_slh__n850), .A (CLOCK_slh__n849));
CLKBUF_X1 CLOCK_slh__c570 (.Z (CLOCK_slh__n851), .A (CLOCK_slh__n850));
CLKBUF_X1 CLOCK_slh__c571 (.Z (CLOCK_slh_n593), .A (CLOCK_slh__n851));
CLKBUF_X1 CLOCK_slh__c575 (.Z (CLOCK_slh__n856), .A (CLOCK_slh__n855));
CLKBUF_X1 CLOCK_slh__c576 (.Z (CLOCK_slh__n857), .A (CLOCK_slh__n856));
CLKBUF_X1 CLOCK_slh__c577 (.Z (CLOCK_slh_n578), .A (CLOCK_slh__n857));
CLKBUF_X1 CLOCK_slh__c581 (.Z (CLOCK_slh__n862), .A (CLOCK_slh__n861));
CLKBUF_X1 CLOCK_slh__c582 (.Z (CLOCK_slh__n863), .A (CLOCK_slh__n862));
CLKBUF_X1 CLOCK_slh__c583 (.Z (CLOCK_slh_n583), .A (CLOCK_slh__n863));
CLKBUF_X1 CLOCK_slh__c587 (.Z (CLOCK_slh__n868), .A (CLOCK_slh__n867));
CLKBUF_X1 CLOCK_slh__c588 (.Z (CLOCK_slh__n869), .A (CLOCK_slh__n868));
CLKBUF_X1 CLOCK_slh__c589 (.Z (CLOCK_slh_n478), .A (CLOCK_slh__n869));
CLKBUF_X1 CLOCK_slh__c593 (.Z (CLOCK_slh__n874), .A (CLOCK_slh__n873));
CLKBUF_X1 CLOCK_slh__c594 (.Z (CLOCK_slh__n875), .A (CLOCK_slh__n874));
CLKBUF_X1 CLOCK_slh__c595 (.Z (CLOCK_slh_n468), .A (CLOCK_slh__n875));
CLKBUF_X1 CLOCK_slh__c599 (.Z (CLOCK_slh__n880), .A (CLOCK_slh__n879));
CLKBUF_X1 CLOCK_slh__c600 (.Z (CLOCK_slh__n881), .A (CLOCK_slh__n880));
CLKBUF_X1 CLOCK_slh__c601 (.Z (CLOCK_slh_n513), .A (CLOCK_slh__n881));
CLKBUF_X1 CLOCK_slh__c605 (.Z (CLOCK_slh__n886), .A (CLOCK_slh__n885));
CLKBUF_X1 CLOCK_slh__c606 (.Z (CLOCK_slh__n887), .A (CLOCK_slh__n886));
CLKBUF_X1 CLOCK_slh__c607 (.Z (CLOCK_slh_n588), .A (CLOCK_slh__n887));
CLKBUF_X1 CLOCK_slh__c611 (.Z (CLOCK_slh__n892), .A (CLOCK_slh__n891));
CLKBUF_X1 CLOCK_slh__c612 (.Z (CLOCK_slh__n893), .A (CLOCK_slh__n892));
CLKBUF_X1 CLOCK_slh__c613 (.Z (CLOCK_slh_n493), .A (CLOCK_slh__n893));
CLKBUF_X1 CLOCK_slh__c617 (.Z (CLOCK_slh__n898), .A (CLOCK_slh__n897));
CLKBUF_X1 CLOCK_slh__c618 (.Z (CLOCK_slh__n899), .A (CLOCK_slh__n898));
CLKBUF_X1 CLOCK_slh__c619 (.Z (CLOCK_slh_n523), .A (CLOCK_slh__n899));
CLKBUF_X1 CLOCK_slh__c623 (.Z (CLOCK_slh__n904), .A (CLOCK_slh__n903));
CLKBUF_X1 CLOCK_slh__c624 (.Z (CLOCK_slh__n905), .A (CLOCK_slh__n904));
CLKBUF_X1 CLOCK_slh__c625 (.Z (CLOCK_slh_n458), .A (CLOCK_slh__n905));
CLKBUF_X1 CLOCK_slh__c629 (.Z (CLOCK_slh__n910), .A (CLOCK_slh__n909));
CLKBUF_X1 CLOCK_slh__c630 (.Z (CLOCK_slh__n911), .A (CLOCK_slh__n910));
CLKBUF_X1 CLOCK_slh__c631 (.Z (CLOCK_slh_n503), .A (CLOCK_slh__n911));
CLKBUF_X1 CLOCK_slh__c635 (.Z (CLOCK_slh__n916), .A (CLOCK_slh__n915));
CLKBUF_X1 CLOCK_slh__c636 (.Z (CLOCK_slh__n917), .A (CLOCK_slh__n916));
CLKBUF_X1 CLOCK_slh__c637 (.Z (CLOCK_slh_n573), .A (CLOCK_slh__n917));
CLKBUF_X1 CLOCK_slh__c641 (.Z (CLOCK_slh__n922), .A (CLOCK_slh__n921));
CLKBUF_X1 CLOCK_slh__c642 (.Z (CLOCK_slh__n923), .A (CLOCK_slh__n922));
CLKBUF_X1 CLOCK_slh__c643 (.Z (CLOCK_slh_n308), .A (CLOCK_slh__n923));
CLKBUF_X1 CLOCK_slh__c647 (.Z (CLOCK_slh__n928), .A (CLOCK_slh__n927));
CLKBUF_X1 CLOCK_slh__c648 (.Z (CLOCK_slh__n929), .A (CLOCK_slh__n928));
CLKBUF_X1 CLOCK_slh__c649 (.Z (CLOCK_slh_n488), .A (CLOCK_slh__n929));
CLKBUF_X1 CLOCK_slh__c653 (.Z (CLOCK_slh__n934), .A (CLOCK_slh__n933));
CLKBUF_X1 CLOCK_slh__c654 (.Z (CLOCK_slh__n935), .A (CLOCK_slh__n934));
CLKBUF_X1 CLOCK_slh__c655 (.Z (CLOCK_slh_n533), .A (CLOCK_slh__n935));
CLKBUF_X1 CLOCK_slh__c659 (.Z (CLOCK_slh__n940), .A (CLOCK_slh__n939));
CLKBUF_X1 CLOCK_slh__c660 (.Z (CLOCK_slh__n941), .A (CLOCK_slh__n940));
CLKBUF_X1 CLOCK_slh__c661 (.Z (CLOCK_slh_n598), .A (CLOCK_slh__n941));
CLKBUF_X1 CLOCK_slh__c665 (.Z (CLOCK_slh__n946), .A (CLOCK_slh__n945));
CLKBUF_X1 CLOCK_slh__c666 (.Z (CLOCK_slh__n947), .A (CLOCK_slh__n946));
CLKBUF_X1 CLOCK_slh__c667 (.Z (CLOCK_slh_n603), .A (CLOCK_slh__n947));
CLKBUF_X1 CLOCK_slh__c671 (.Z (CLOCK_slh__n952), .A (CLOCK_slh__n951));
CLKBUF_X1 CLOCK_slh__c672 (.Z (CLOCK_slh__n953), .A (CLOCK_slh__n952));
CLKBUF_X1 CLOCK_slh__c673 (.Z (CLOCK_slh_n608), .A (CLOCK_slh__n953));
CLKBUF_X1 CLOCK_slh__c677 (.Z (CLOCK_slh__n958), .A (CLOCK_slh__n957));
CLKBUF_X1 CLOCK_slh__c678 (.Z (CLOCK_slh__n959), .A (CLOCK_slh__n958));
CLKBUF_X1 CLOCK_slh__c679 (.Z (CLOCK_slh_n618), .A (CLOCK_slh__n959));
CLKBUF_X1 CLOCK_slh__c683 (.Z (CLOCK_slh__n964), .A (CLOCK_slh__n963));
CLKBUF_X1 CLOCK_slh__c684 (.Z (CLOCK_slh__n965), .A (CLOCK_slh__n964));
CLKBUF_X1 CLOCK_slh__c685 (.Z (CLOCK_slh_n553), .A (CLOCK_slh__n965));
CLKBUF_X1 CLOCK_slh__c689 (.Z (CLOCK_slh__n970), .A (CLOCK_slh__n969));
CLKBUF_X1 CLOCK_slh__c690 (.Z (CLOCK_slh__n971), .A (CLOCK_slh__n970));
CLKBUF_X1 CLOCK_slh__c691 (.Z (CLOCK_slh_n453), .A (CLOCK_slh__n971));
CLKBUF_X1 CLOCK_slh__c695 (.Z (CLOCK_slh__n976), .A (CLOCK_slh__n975));
CLKBUF_X1 CLOCK_slh__c696 (.Z (CLOCK_slh__n977), .A (CLOCK_slh__n976));
CLKBUF_X1 CLOCK_slh__c697 (.Z (CLOCK_slh_n323), .A (CLOCK_slh__n977));
CLKBUF_X1 CLOCK_slh__c701 (.Z (CLOCK_slh__n982), .A (CLOCK_slh__n981));
CLKBUF_X1 CLOCK_slh__c702 (.Z (CLOCK_slh__n983), .A (CLOCK_slh__n982));
CLKBUF_X1 CLOCK_slh__c703 (.Z (CLOCK_slh_n443), .A (CLOCK_slh__n983));
CLKBUF_X1 CLOCK_slh__c707 (.Z (CLOCK_slh__n988), .A (CLOCK_slh__n987));
CLKBUF_X1 CLOCK_slh__c708 (.Z (CLOCK_slh__n989), .A (CLOCK_slh__n988));
CLKBUF_X1 CLOCK_slh__c709 (.Z (CLOCK_slh_n613), .A (CLOCK_slh__n989));
CLKBUF_X1 CLOCK_slh__c713 (.Z (CLOCK_slh__n994), .A (CLOCK_slh__n993));
CLKBUF_X1 CLOCK_slh__c714 (.Z (CLOCK_slh__n995), .A (CLOCK_slh__n994));
CLKBUF_X1 CLOCK_slh__c715 (.Z (CLOCK_slh_n428), .A (CLOCK_slh__n995));
CLKBUF_X1 CLOCK_slh__c719 (.Z (CLOCK_slh__n1000), .A (CLOCK_slh__n999));
CLKBUF_X1 CLOCK_slh__c720 (.Z (CLOCK_slh__n1001), .A (CLOCK_slh__n1000));
CLKBUF_X1 CLOCK_slh__c721 (.Z (CLOCK_slh_n313), .A (CLOCK_slh__n1001));
CLKBUF_X1 CLOCK_slh__c725 (.Z (CLOCK_slh__n1006), .A (CLOCK_slh__n1005));
CLKBUF_X1 CLOCK_slh__c726 (.Z (CLOCK_slh__n1007), .A (CLOCK_slh__n1006));
CLKBUF_X1 CLOCK_slh__c727 (.Z (CLOCK_slh_n543), .A (CLOCK_slh__n1007));
CLKBUF_X1 CLOCK_slh__c731 (.Z (CLOCK_slh__n1012), .A (CLOCK_slh__n1011));
CLKBUF_X1 CLOCK_slh__c732 (.Z (CLOCK_slh__n1013), .A (CLOCK_slh__n1012));
CLKBUF_X1 CLOCK_slh__c733 (.Z (CLOCK_slh_n368), .A (CLOCK_slh__n1013));
CLKBUF_X1 CLOCK_slh__c737 (.Z (CLOCK_slh__n1018), .A (CLOCK_slh__n1017));
CLKBUF_X1 CLOCK_slh__c738 (.Z (CLOCK_slh__n1019), .A (CLOCK_slh__n1018));
CLKBUF_X1 CLOCK_slh__c739 (.Z (CLOCK_slh_n433), .A (CLOCK_slh__n1019));

endmodule //Radix4


