
// 	Fri Dec 23 04:16:03 2022
//	vlsi
//	localhost.localdomain

module registerNbits (clk_CTS_1_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_3;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_2), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_2), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_2), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid0_2), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid0_2), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid0_2), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_2), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid0_2), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid0_2), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid0_2), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid0_2), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid0_2), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid0_2), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_2), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_2), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_2), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_2), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_2), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_2), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_2), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_2), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_2), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_2), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_2), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_2), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_2), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_2), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_2), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_2), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_2), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_2), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid0_2), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid0_3), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L3_c_tid0_3 (.Z (CTS_n_tid0_2), .A (CTS_n_tid0_3));

endmodule //registerNbits

module registerNbits__2_8 (clk_CTS_1_PP_0, clk_CTS_1_PP_1, clk, reset, en, inp, out);

output [31:0] out;
output clk_CTS_1_PP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_1;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_3;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_2), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_2), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_2), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_2), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_2), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_2), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_2), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_2), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_2), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_2), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_2), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_2), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_2), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_2), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_2), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_2), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_2), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_2), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_2), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_2), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_2), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_2), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_2), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_2), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_2), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_2), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_2), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_2), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_2), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_2), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_2), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_2), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid1_3), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L3_c_tid1_3 (.Z (CTS_n_tid1_2), .A (CTS_n_tid1_3));
CLKBUF_X3 CTS_L1_c_tid1_42 (.Z (clk_CTS_1_PP_0), .A (clk_CTS_1_PP_1));

endmodule //registerNbits__2_8

module registerNbits__2_5 (clk_CTS_1_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_0;
wire drc_ipo_n180;
wire drc_ipo_n178;
wire drc_ipo_n176;
wire drc_ipo_n174;
wire drc_ipo_n172;
wire drc_ipo_n170;
wire drc_ipo_n168;
wire drc_ipo_n166;
wire drc_ipo_n164;
wire drc_ipo_n162;
wire drc_ipo_n160;
wire drc_ipo_n158;
wire drc_ipo_n156;
wire drc_ipo_n154;
wire drc_ipo_n152;
wire drc_ipo_n150;
wire drc_ipo_n148;
wire drc_ipo_n146;
wire drc_ipo_n144;
wire drc_ipo_n142;
wire drc_ipo_n140;
wire drc_ipo_n138;
wire drc_ipo_n136;
wire drc_ipo_n134;
wire drc_ipo_n132;
wire drc_ipo_n130;
wire drc_ipo_n128;
wire drc_ipo_n126;
wire drc_ipo_n124;
wire drc_ipo_n122;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_182;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_183;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_182), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_182), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (drc_ipo_n122), .CK (CTS_n_tid0_182), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (drc_ipo_n124), .CK (CTS_n_tid0_182), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (drc_ipo_n126), .CK (CTS_n_tid0_182), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (drc_ipo_n128), .CK (CTS_n_tid0_182), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (drc_ipo_n130), .CK (CTS_n_tid0_182), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (drc_ipo_n132), .CK (CTS_n_tid0_182), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (drc_ipo_n134), .CK (CTS_n_tid0_182), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (drc_ipo_n136), .CK (CTS_n_tid0_182), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (drc_ipo_n138), .CK (CTS_n_tid0_182), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (drc_ipo_n140), .CK (CTS_n_tid0_182), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (drc_ipo_n142), .CK (CTS_n_tid0_182), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (drc_ipo_n144), .CK (CTS_n_tid0_182), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (drc_ipo_n146), .CK (CTS_n_tid0_182), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (drc_ipo_n148), .CK (CTS_n_tid0_182), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (drc_ipo_n150), .CK (CTS_n_tid0_182), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (drc_ipo_n152), .CK (CTS_n_tid0_182), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (drc_ipo_n154), .CK (CTS_n_tid0_182), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (drc_ipo_n156), .CK (CTS_n_tid0_182), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (drc_ipo_n158), .CK (CTS_n_tid0_182), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (drc_ipo_n160), .CK (CTS_n_tid0_182), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (drc_ipo_n162), .CK (CTS_n_tid0_182), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (drc_ipo_n164), .CK (CTS_n_tid0_182), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (drc_ipo_n166), .CK (CTS_n_tid0_182), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (drc_ipo_n168), .CK (CTS_n_tid0_182), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (drc_ipo_n170), .CK (CTS_n_tid0_182), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (drc_ipo_n172), .CK (CTS_n_tid0_182), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (drc_ipo_n174), .CK (CTS_n_tid0_182), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (drc_ipo_n176), .CK (CTS_n_tid0_182), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (drc_ipo_n178), .CK (CTS_n_tid0_182), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n180), .CK (CTS_n_tid0_182), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid0_183), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X2 drc_ipo_c90 (.Z (out[31]), .A (drc_ipo_n180));
CLKBUF_X2 drc_ipo_c89 (.Z (out[30]), .A (drc_ipo_n178));
CLKBUF_X2 drc_ipo_c88 (.Z (out[29]), .A (drc_ipo_n176));
CLKBUF_X2 drc_ipo_c87 (.Z (out[28]), .A (drc_ipo_n174));
CLKBUF_X2 drc_ipo_c86 (.Z (out[27]), .A (drc_ipo_n172));
CLKBUF_X2 drc_ipo_c85 (.Z (out[26]), .A (drc_ipo_n170));
CLKBUF_X2 drc_ipo_c84 (.Z (out[25]), .A (drc_ipo_n168));
CLKBUF_X2 drc_ipo_c83 (.Z (out[24]), .A (drc_ipo_n166));
CLKBUF_X2 drc_ipo_c82 (.Z (out[23]), .A (drc_ipo_n164));
CLKBUF_X2 drc_ipo_c81 (.Z (out[22]), .A (drc_ipo_n162));
CLKBUF_X2 drc_ipo_c80 (.Z (out[21]), .A (drc_ipo_n160));
CLKBUF_X2 drc_ipo_c79 (.Z (out[20]), .A (drc_ipo_n158));
CLKBUF_X2 drc_ipo_c78 (.Z (out[19]), .A (drc_ipo_n156));
CLKBUF_X2 drc_ipo_c77 (.Z (out[18]), .A (drc_ipo_n154));
CLKBUF_X2 drc_ipo_c76 (.Z (out[17]), .A (drc_ipo_n152));
CLKBUF_X2 drc_ipo_c75 (.Z (out[16]), .A (drc_ipo_n150));
CLKBUF_X2 drc_ipo_c74 (.Z (out[15]), .A (drc_ipo_n148));
CLKBUF_X2 drc_ipo_c73 (.Z (out[14]), .A (drc_ipo_n146));
CLKBUF_X2 drc_ipo_c72 (.Z (out[13]), .A (drc_ipo_n144));
CLKBUF_X2 drc_ipo_c71 (.Z (out[12]), .A (drc_ipo_n142));
BUF_X4 drc_ipo_c70 (.Z (out[11]), .A (drc_ipo_n140));
CLKBUF_X2 drc_ipo_c69 (.Z (out[10]), .A (drc_ipo_n138));
CLKBUF_X2 drc_ipo_c68 (.Z (out[9]), .A (drc_ipo_n136));
CLKBUF_X2 drc_ipo_c67 (.Z (out[8]), .A (drc_ipo_n134));
CLKBUF_X2 drc_ipo_c66 (.Z (out[7]), .A (drc_ipo_n132));
CLKBUF_X2 drc_ipo_c65 (.Z (out[6]), .A (drc_ipo_n130));
CLKBUF_X2 drc_ipo_c64 (.Z (out[5]), .A (drc_ipo_n128));
CLKBUF_X2 drc_ipo_c63 (.Z (out[4]), .A (drc_ipo_n126));
CLKBUF_X2 drc_ipo_c62 (.Z (out[3]), .A (drc_ipo_n124));
CLKBUF_X2 drc_ipo_c61 (.Z (out[2]), .A (drc_ipo_n122));
CLKBUF_X3 CTS_L3_c_tid0_93 (.Z (CTS_n_tid0_182), .A (CTS_n_tid0_183));

endmodule //registerNbits__2_5

module registerNbits__2_2 (clk_CTS_1_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_0;
wire drc_ipo_n186;
wire drc_ipo_n184;
wire drc_ipo_n182;
wire drc_ipo_n180;
wire drc_ipo_n178;
wire drc_ipo_n176;
wire drc_ipo_n174;
wire drc_ipo_n172;
wire drc_ipo_n170;
wire drc_ipo_n168;
wire drc_ipo_n166;
wire drc_ipo_n164;
wire drc_ipo_n162;
wire drc_ipo_n160;
wire drc_ipo_n158;
wire drc_ipo_n156;
wire drc_ipo_n154;
wire drc_ipo_n152;
wire drc_ipo_n150;
wire drc_ipo_n148;
wire drc_ipo_n146;
wire drc_ipo_n144;
wire drc_ipo_n142;
wire drc_ipo_n140;
wire drc_ipo_n138;
wire drc_ipo_n136;
wire drc_ipo_n134;
wire drc_ipo_n132;
wire drc_ipo_n130;
wire drc_ipo_n128;
wire drc_ipo_n126;
wire n_0_0;
wire n_1;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_192;
wire CTS_n_tid1_193;
wire CTS_n_tid1_194;
wire CTS_n_tid1_195;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (drc_ipo_n126), .CK (CTS_n_tid1_194), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (drc_ipo_n128), .CK (CTS_n_tid1_193), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (drc_ipo_n130), .CK (CTS_n_tid1_193), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (drc_ipo_n132), .CK (CTS_n_tid1_193), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (drc_ipo_n134), .CK (CTS_n_tid1_193), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (drc_ipo_n136), .CK (CTS_n_tid1_193), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (drc_ipo_n138), .CK (CTS_n_tid1_193), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (drc_ipo_n140), .CK (CTS_n_tid1_193), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (drc_ipo_n142), .CK (CTS_n_tid1_194), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (drc_ipo_n144), .CK (CTS_n_tid1_195), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (drc_ipo_n146), .CK (CTS_n_tid1_193), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (drc_ipo_n148), .CK (CTS_n_tid1_195), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (drc_ipo_n150), .CK (CTS_n_tid1_195), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (drc_ipo_n152), .CK (CTS_n_tid1_195), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (drc_ipo_n154), .CK (CTS_n_tid1_194), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (drc_ipo_n156), .CK (CTS_n_tid1_194), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (drc_ipo_n158), .CK (CTS_n_tid1_195), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (drc_ipo_n160), .CK (CTS_n_tid1_195), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (drc_ipo_n162), .CK (CTS_n_tid1_195), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (drc_ipo_n164), .CK (CTS_n_tid1_194), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (drc_ipo_n166), .CK (CTS_n_tid1_194), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (drc_ipo_n168), .CK (CTS_n_tid1_195), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (drc_ipo_n170), .CK (CTS_n_tid1_195), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (drc_ipo_n172), .CK (CTS_n_tid1_194), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (drc_ipo_n174), .CK (CTS_n_tid1_195), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (drc_ipo_n176), .CK (CTS_n_tid1_194), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (drc_ipo_n178), .CK (CTS_n_tid1_194), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (drc_ipo_n180), .CK (CTS_n_tid1_195), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (drc_ipo_n182), .CK (CTS_n_tid1_194), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (drc_ipo_n184), .CK (CTS_n_tid1_194), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_194), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n186), .CK (CTS_n_tid1_194), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid1_192), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X2 drc_ipo_c93 (.Z (out[31]), .A (drc_ipo_n186));
CLKBUF_X2 drc_ipo_c92 (.Z (out[29]), .A (drc_ipo_n184));
CLKBUF_X2 drc_ipo_c91 (.Z (out[28]), .A (drc_ipo_n182));
CLKBUF_X2 drc_ipo_c90 (.Z (out[27]), .A (drc_ipo_n180));
CLKBUF_X2 drc_ipo_c89 (.Z (out[26]), .A (drc_ipo_n178));
CLKBUF_X2 drc_ipo_c88 (.Z (out[25]), .A (drc_ipo_n176));
CLKBUF_X2 drc_ipo_c87 (.Z (out[24]), .A (drc_ipo_n174));
CLKBUF_X2 drc_ipo_c86 (.Z (out[23]), .A (drc_ipo_n172));
CLKBUF_X2 drc_ipo_c85 (.Z (out[22]), .A (drc_ipo_n170));
CLKBUF_X2 drc_ipo_c84 (.Z (out[21]), .A (drc_ipo_n168));
CLKBUF_X2 drc_ipo_c83 (.Z (out[20]), .A (drc_ipo_n166));
CLKBUF_X2 drc_ipo_c82 (.Z (out[19]), .A (drc_ipo_n164));
CLKBUF_X2 drc_ipo_c81 (.Z (out[18]), .A (drc_ipo_n162));
CLKBUF_X2 drc_ipo_c80 (.Z (out[17]), .A (drc_ipo_n160));
CLKBUF_X2 drc_ipo_c79 (.Z (out[16]), .A (drc_ipo_n158));
CLKBUF_X2 drc_ipo_c78 (.Z (out[15]), .A (drc_ipo_n156));
CLKBUF_X2 drc_ipo_c77 (.Z (out[14]), .A (drc_ipo_n154));
CLKBUF_X2 drc_ipo_c76 (.Z (out[13]), .A (drc_ipo_n152));
CLKBUF_X2 drc_ipo_c75 (.Z (out[12]), .A (drc_ipo_n150));
CLKBUF_X2 drc_ipo_c74 (.Z (out[11]), .A (drc_ipo_n148));
BUF_X4 drc_ipo_c73 (.Z (out[10]), .A (drc_ipo_n146));
CLKBUF_X2 drc_ipo_c72 (.Z (out[9]), .A (drc_ipo_n144));
CLKBUF_X2 drc_ipo_c71 (.Z (out[8]), .A (drc_ipo_n142));
CLKBUF_X2 drc_ipo_c70 (.Z (out[7]), .A (drc_ipo_n140));
CLKBUF_X2 drc_ipo_c69 (.Z (out[6]), .A (drc_ipo_n138));
CLKBUF_X2 drc_ipo_c68 (.Z (out[5]), .A (drc_ipo_n136));
CLKBUF_X2 drc_ipo_c67 (.Z (out[4]), .A (drc_ipo_n134));
CLKBUF_X2 drc_ipo_c66 (.Z (out[3]), .A (drc_ipo_n132));
CLKBUF_X2 drc_ipo_c65 (.Z (out[2]), .A (drc_ipo_n130));
CLKBUF_X2 drc_ipo_c64 (.Z (out[1]), .A (drc_ipo_n128));
CLKBUF_X2 drc_ipo_c63 (.Z (out[0]), .A (drc_ipo_n126));
CLKBUF_X3 CTS_L3_c_tid1_98 (.Z (CTS_n_tid1_193), .A (CTS_n_tid1_192));
CLKBUF_X3 CTS_L3_c_tid1_99 (.Z (CTS_n_tid1_194), .A (CTS_n_tid1_192));
CLKBUF_X3 CTS_L3_c_tid1_100 (.Z (CTS_n_tid1_195), .A (CTS_n_tid1_192));

endmodule //registerNbits__2_2

module datapath (inputB, inputA, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;
wire n_3;
wire n_51;
wire n_2366;
wire n_2371;
wire n_2367;
wire n_36;
wire n_9;
wire n_61;
wire n_10;
wire n_11;
wire n_2363;
wire n_2362;
wire n_42;
wire n_43;
wire n_72;
wire n_44;
wire n_73;
wire n_78;
wire n_45;
wire n_46;
wire n_12;
wire n_2364;
wire n_2365;
wire n_55;
wire n_13;
wire n_2359;
wire n_2357;
wire n_64;
wire n_65;
wire n_2379;
wire n_2375;
wire n_90;
wire n_2355;
wire n_2356;
wire n_93;
wire n_94;
wire n_95;
wire n_2373;
wire n_2374;
wire n_2380;
wire n_108;
wire n_2350;
wire n_119;
wire n_120;
wire n_121;
wire n_2381;
wire n_134;
wire n_2337;
wire n_2349;
wire n_2338;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_2336;
wire n_2372;
wire n_166;
wire n_2331;
wire n_2321;
wire n_197;
wire n_198;
wire n_199;
wire n_2327;
wire n_2325;
wire n_2329;
wire n_2328;
wire n_220;
wire n_2233;
wire n_2214;
wire n_229;
wire n_231;
wire n_2195;
wire n_232;
wire n_2241;
wire n_233;
wire n_234;
wire n_235;
wire n_2259;
wire n_236;
wire n_2319;
wire n_2335;
wire n_2320;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_2291;
wire n_2287;
wire n_2292;
wire n_2312;
wire n_244;
wire n_2289;
wire n_2288;
wire n_2290;
wire n_2203;
wire n_245;
wire n_2314;
wire n_690;
wire n_1349;
wire n_2186;
wire n_1219;
wire n_864;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_2246;
wire n_2204;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_2260;
wire n_2286;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_2187;
wire n_306;
wire n_14;
wire n_2433;
wire n_2434;
wire n_2529;
wire n_320;
wire n_2170;
wire n_321;
wire n_322;
wire n_323;
wire n_2208;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_324;
wire n_2249;
wire n_2248;
wire n_2247;
wire n_325;
wire n_326;
wire n_15;
wire n_2439;
wire n_2140;
wire n_332;
wire n_335;
wire n_2422;
wire n_336;
wire n_337;
wire n_2451;
wire n_2441;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_2188;
wire n_2196;
wire n_357;
wire n_2436;
wire n_2432;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_2423;
wire n_2420;
wire n_374;
wire n_2421;
wire n_377;
wire n_2182;
wire n_378;
wire n_2171;
wire n_2174;
wire n_379;
wire n_380;
wire n_2131;
wire n_2130;
wire n_386;
wire n_387;
wire n_2430;
wire n_2429;
wire n_391;
wire n_2122;
wire n_2121;
wire n_396;
wire n_2137;
wire n_2136;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_16;
wire n_2501;
wire n_2489;
wire n_434;
wire n_435;
wire n_2506;
wire n_2502;
wire n_453;
wire n_454;
wire n_455;
wire n_2424;
wire n_2418;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_2484;
wire n_2483;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_2110;
wire n_2119;
wire n_519;
wire n_520;
wire n_2415;
wire n_2414;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_2524;
wire n_2482;
wire n_580;
wire n_2413;
wire n_2453;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_2411;
wire n_2478;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_2412;
wire n_695;
wire n_2456;
wire n_2458;
wire n_2457;
wire n_696;
wire n_1806;
wire n_1801;
wire n_713;
wire n_1992;
wire n_1991;
wire n_718;
wire n_1988;
wire n_1987;
wire n_724;
wire n_725;
wire n_1980;
wire n_1978;
wire n_732;
wire n_733;
wire n_734;
wire n_2475;
wire n_2459;
wire n_2477;
wire n_2476;
wire n_735;
wire n_736;
wire n_737;
wire n_2083;
wire n_2038;
wire n_771;
wire n_772;
wire n_2410;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_2059;
wire n_2077;
wire n_2082;
wire n_2078;
wire n_782;
wire n_783;
wire n_1983;
wire n_1976;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_1797;
wire n_1796;
wire n_817;
wire n_818;
wire n_2057;
wire n_819;
wire n_2039;
wire n_2056;
wire n_2058;
wire n_820;
wire n_2006;
wire n_2004;
wire n_840;
wire n_1998;
wire n_2000;
wire n_1999;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_2037;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_1931;
wire n_1930;
wire n_926;
wire n_927;
wire n_928;
wire n_930;
wire n_931;
wire n_1795;
wire n_932;
wire n_933;
wire n_934;
wire n_2558;
wire n_945;
wire n_2557;
wire n_947;
wire n_2564;
wire n_955;
wire n_956;
wire n_1794;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_1965;
wire n_1932;
wire n_974;
wire n_975;
wire n_976;
wire n_1901;
wire n_977;
wire n_1902;
wire n_1903;
wire n_1896;
wire n_978;
wire n_2555;
wire n_2552;
wire n_1723;
wire n_2551;
wire n_979;
wire n_2560;
wire n_2562;
wire n_2563;
wire n_980;
wire n_981;
wire n_982;
wire n_2656;
wire n_984;
wire n_985;
wire n_986;
wire n_1724;
wire n_400;
wire n_987;
wire n_988;
wire n_2740;
wire n_990;
wire n_991;
wire n_992;
wire n_2559;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_2622;
wire n_2615;
wire n_1013;
wire n_1014;
wire n_2587;
wire n_2585;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_2578;
wire n_2581;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_2566;
wire n_2577;
wire n_2574;
wire n_2576;
wire n_1074;
wire n_2583;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_2550;
wire n_2565;
wire n_2543;
wire n_2549;
wire n_1092;
wire n_2692;
wire n_2685;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_67;
wire n_414;
wire n_1110;
wire n_1111;
wire n_66;
wire n_217;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_2633;
wire n_2630;
wire n_2629;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_2651;
wire n_2650;
wire n_1125;
wire n_1128;
wire n_2647;
wire n_1129;
wire n_1130;
wire n_1133;
wire n_2654;
wire n_1134;
wire n_1135;
wire n_2679;
wire n_2681;
wire n_2680;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_2582;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_2607;
wire n_1174;
wire n_2606;
wire n_2604;
wire n_2612;
wire n_1175;
wire n_1176;
wire n_2675;
wire n_1177;
wire n_1178;
wire n_2635;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_2880;
wire n_2879;
wire n_1218;
wire n_2894;
wire n_2884;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_2613;
wire n_1236;
wire n_2584;
wire n_2602;
wire n_2603;
wire n_1237;
wire n_2751;
wire n_2750;
wire n_1242;
wire n_2746;
wire n_2745;
wire n_1248;
wire n_1249;
wire n_2717;
wire n_2764;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_2636;
wire n_2657;
wire n_1279;
wire n_2800;
wire n_2799;
wire n_1299;
wire n_2794;
wire n_2793;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_2760;
wire n_2759;
wire n_1328;
wire n_1329;
wire n_2741;
wire n_2715;
wire n_1335;
wire n_1336;
wire n_2676;
wire n_1337;
wire n_1338;
wire n_2903;
wire n_2873;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_2771;
wire n_2765;
wire n_1362;
wire n_2902;
wire n_2900;
wire n_2899;
wire n_1363;
wire n_2890;
wire n_2888;
wire n_2887;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_2755;
wire n_2754;
wire n_1397;
wire n_2714;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1437;
wire n_1438;
wire n_3543;
wire n_2959;
wire n_1444;
wire n_3538;
wire n_3537;
wire n_1448;
wire n_1449;
wire n_3510;
wire n_3509;
wire n_1454;
wire n_1455;
wire n_2850;
wire n_3047;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_3071;
wire n_1461;
wire n_3517;
wire n_3518;
wire n_3534;
wire n_1468;
wire n_1469;
wire n_3215;
wire n_3214;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_2924;
wire n_2923;
wire n_2926;
wire n_2925;
wire n_1479;
wire n_3007;
wire n_1481;
wire n_63;
wire n_585;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1490;
wire n_3562;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_2789;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_2804;
wire n_2791;
wire n_2792;
wire n_2798;
wire n_1505;
wire n_2815;
wire n_1506;
wire n_2814;
wire n_2809;
wire n_2819;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_2979;
wire n_2978;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_2825;
wire n_2808;
wire n_2831;
wire n_2826;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_2806;
wire n_2790;
wire n_2851;
wire n_2807;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1539;
wire n_17;
wire n_3507;
wire n_1541;
wire n_3540;
wire n_3536;
wire n_1548;
wire n_1549;
wire n_3218;
wire n_3206;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_2941;
wire n_2940;
wire n_1578;
wire n_3048;
wire n_1583;
wire n_1584;
wire n_1587;
wire n_3040;
wire n_1588;
wire n_1589;
wire n_2697;
wire n_1590;
wire n_2964;
wire n_2963;
wire n_1596;
wire n_2955;
wire n_2954;
wire n_1601;
wire n_1602;
wire n_2950;
wire n_2949;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_3500;
wire n_3499;
wire n_1654;
wire n_1655;
wire n_2712;
wire n_2698;
wire n_2706;
wire n_2700;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_3535;
wire n_3480;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_2934;
wire n_2933;
wire n_1683;
wire n_1686;
wire n_3381;
wire n_1687;
wire n_2968;
wire n_1688;
wire n_18;
wire n_1690;
wire n_1691;
wire n_3377;
wire n_3376;
wire n_1695;
wire n_1696;
wire n_19;
wire n_20;
wire n_21;
wire n_3489;
wire n_3491;
wire n_3490;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_3200;
wire n_3199;
wire n_1734;
wire n_2970;
wire n_2961;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1774;
wire n_2927;
wire n_1775;
wire n_1776;
wire n_22;
wire n_3182;
wire n_3195;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_3496;
wire n_3488;
wire n_1830;
wire n_3316;
wire n_3315;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_3477;
wire n_3475;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_3179;
wire n_3072;
wire n_1906;
wire n_3485;
wire n_3473;
wire n_1920;
wire n_1921;
wire n_1604;
wire n_23;
wire n_1515;
wire n_24;
wire n_1605;
wire n_25;
wire n_1941;
wire n_1942;
wire n_3008;
wire n_1943;
wire n_3312;
wire n_3320;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_3168;
wire n_1471;
wire n_26;
wire n_27;
wire n_3247;
wire n_3246;
wire n_1977;
wire n_4162;
wire n_314;
wire n_1136;
wire n_1979;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_3418;
wire n_3417;
wire n_1996;
wire n_1997;
wire n_3256;
wire n_3268;
wire n_3273;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_3464;
wire n_3463;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_3138;
wire n_32;
wire n_3469;
wire n_3468;
wire n_2123;
wire n_3253;
wire n_33;
wire n_3353;
wire n_3349;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_3323;
wire n_3301;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_3467;
wire n_3459;
wire n_2177;
wire n_3233;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_853;
wire n_34;
wire n_35;
wire n_3300;
wire n_3297;
wire n_2256;
wire n_529;
wire n_530;
wire n_881;
wire n_37;
wire n_38;
wire n_3348;
wire n_3327;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_39;
wire n_1661;
wire n_1660;
wire n_2332;
wire n_3235;
wire n_3234;
wire n_3291;
wire n_3236;
wire n_2333;
wire n_2334;
wire n_1719;
wire n_1718;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_833;
wire n_40;
wire n_1514;
wire n_41;
wire n_3455;
wire n_3454;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_1711;
wire n_1653;
wire n_2474;
wire n_895;
wire n_893;
wire n_2490;
wire n_47;
wire n_1146;
wire n_1148;
wire n_1147;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_1143;
wire n_1142;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_1559;
wire n_1554;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2575;
wire n_3294;
wire n_2591;
wire n_3453;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_1649;
wire n_1553;
wire n_2614;
wire n_899;
wire n_892;
wire n_2631;
wire n_1139;
wire n_1152;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_1312;
wire n_1225;
wire n_2663;
wire n_701;
wire n_702;
wire n_2682;
wire n_680;
wire n_681;
wire n_2699;
wire n_674;
wire n_675;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_3408;
wire n_2723;
wire n_3295;
wire n_3400;
wire n_3407;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2778;
wire n_1350;
wire n_2779;
wire n_1552;
wire n_2780;
wire n_2781;
wire n_1222;
wire n_1221;
wire n_2827;
wire n_703;
wire n_707;
wire n_2832;
wire n_648;
wire n_590;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_4109;
wire n_756;
wire n_2878;
wire n_2881;
wire n_4133;
wire n_48;
wire n_1016;
wire n_49;
wire n_4135;
wire n_2885;
wire n_2886;
wire n_4129;
wire n_4128;
wire n_2892;
wire n_2893;
wire n_4119;
wire n_4118;
wire n_2897;
wire n_50;
wire n_4159;
wire n_4160;
wire n_4163;
wire n_2905;
wire n_2906;
wire n_4150;
wire n_4149;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_1137;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_1220;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_1361;
wire n_2972;
wire n_1355;
wire n_1357;
wire n_1359;
wire n_2973;
wire n_710;
wire n_2974;
wire n_2981;
wire n_4157;
wire n_2982;
wire n_2983;
wire n_767;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_763;
wire n_4060;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_1551;
wire n_127;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_709;
wire n_2997;
wire n_589;
wire n_2999;
wire n_3000;
wire n_883;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_940;
wire n_884;
wire n_1017;
wire n_942;
wire n_3005;
wire n_719;
wire n_714;
wire n_715;
wire n_717;
wire n_3006;
wire n_4062;
wire n_3010;
wire n_4058;
wire n_4057;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_4345;
wire n_4344;
wire n_3021;
wire n_4319;
wire n_4028;
wire n_3027;
wire n_3028;
wire n_4051;
wire n_4050;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_4353;
wire n_4351;
wire n_3041;
wire n_3044;
wire n_4367;
wire n_3045;
wire n_3046;
wire n_4335;
wire n_4334;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_1049;
wire n_3066;
wire n_1038;
wire n_1019;
wire n_1039;
wire n_3067;
wire n_1020;
wire n_1029;
wire n_1021;
wire n_1024;
wire n_3068;
wire n_1006;
wire n_1005;
wire n_999;
wire n_3069;
wire n_3070;
wire n_4099;
wire n_4098;
wire n_3076;
wire n_3077;
wire n_943;
wire n_3078;
wire n_952;
wire n_3079;
wire n_951;
wire n_998;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_757;
wire n_3086;
wire n_721;
wire n_3087;
wire n_720;
wire n_711;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_4154;
wire n_4136;
wire n_3100;
wire n_4123;
wire n_4117;
wire n_3108;
wire n_3109;
wire n_1040;
wire n_3110;
wire n_1041;
wire n_1048;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_4082;
wire n_4067;
wire n_3135;
wire n_3139;
wire n_4065;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3961;
wire n_3960;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3988;
wire n_3987;
wire n_3173;
wire n_3980;
wire n_3979;
wire n_3180;
wire n_3181;
wire n_3971;
wire n_3970;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_4364;
wire n_4350;
wire n_3197;
wire n_4061;
wire n_4042;
wire n_3202;
wire n_3203;
wire n_4321;
wire n_4316;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_4112;
wire n_4097;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_4312;
wire n_4311;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3965;
wire n_3959;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_4086;
wire n_4035;
wire n_3282;
wire n_4301;
wire n_4303;
wire n_4302;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3681;
wire n_3680;
wire n_3317;
wire n_3716;
wire n_3715;
wire n_3321;
wire n_3322;
wire n_3672;
wire n_3671;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_4034;
wire n_3945;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_4197;
wire n_4196;
wire n_3375;
wire n_4234;
wire n_4233;
wire n_3379;
wire n_3380;
wire n_4242;
wire n_4241;
wire n_3384;
wire n_3385;
wire n_3388;
wire n_4259;
wire n_3389;
wire n_4261;
wire n_3788;
wire n_3395;
wire n_3396;
wire n_4248;
wire n_3689;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_4296;
wire n_4291;
wire n_3419;
wire n_3677;
wire n_3670;
wire n_3427;
wire n_4175;
wire n_4169;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_4290;
wire n_4276;
wire n_3494;
wire n_3495;
wire n_4256;
wire n_4245;
wire n_3502;
wire n_4295;
wire n_3503;
wire n_4293;
wire n_4292;
wire n_4294;
wire n_3504;
wire n_3505;
wire n_3642;
wire n_3628;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_4238;
wire n_4232;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3944;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_4192;
wire n_4168;
wire n_3546;
wire n_3948;
wire n_3547;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3573;
wire n_3574;
wire n_4164;
wire n_3575;
wire n_4275;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3891;
wire n_3890;
wire n_3599;
wire n_3600;
wire n_3907;
wire n_3897;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3721;
wire n_3627;
wire n_3633;
wire n_3634;
wire n_4279;
wire n_4285;
wire n_4280;
wire n_4282;
wire n_3635;
wire n_3821;
wire n_3801;
wire n_3643;
wire n_3644;
wire n_4287;
wire n_4286;
wire n_4289;
wire n_4288;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_578;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_584;
wire n_3688;
wire n_3624;
wire n_577;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_588;
wire n_215;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_213;
wire n_3696;
wire n_216;
wire n_259;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3789;
wire n_3704;
wire n_3705;
wire n_4218;
wire n_4165;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_4244;
wire n_4220;
wire n_4227;
wire n_4221;
wire n_3714;
wire n_3588;
wire n_3572;
wire n_3719;
wire n_3720;
wire n_3610;
wire n_3605;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3626;
wire n_3732;
wire n_3568;
wire n_3567;
wire n_3738;
wire n_3740;
wire n_510;
wire n_3741;
wire n_3596;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3602;
wire n_513;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_478;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_493;
wire n_492;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_512;
wire n_511;
wire n_3792;
wire n_567;
wire n_566;
wire n_3798;
wire n_506;
wire n_500;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3564;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3790;
wire n_3888;
wire n_3896;
wire n_3889;
wire n_3813;
wire n_3794;
wire n_3793;
wire n_3795;
wire n_3815;
wire n_3818;
wire n_575;
wire n_3819;
wire n_579;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3799;
wire n_3791;
wire n_3871;
wire n_3800;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3604;
wire n_3565;
wire n_3571;
wire n_3566;
wire n_3851;
wire n_515;
wire n_514;
wire n_3857;
wire n_522;
wire n_521;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_482;
wire n_461;
wire n_218;
wire n_3868;
wire n_3869;
wire n_509;
wire n_3870;
wire n_570;
wire n_389;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_583;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_571;
wire n_565;
wire n_3893;
wire n_495;
wire n_491;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_556;
wire n_574;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_442;
wire n_443;
wire n_445;
wire n_3942;
wire n_3943;
wire n_490;
wire n_486;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_561;
wire n_559;
wire n_3968;
wire n_551;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_546;
wire n_544;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_282;
wire n_281;
wire n_4011;
wire n_4012;
wire n_555;
wire n_4013;
wire n_553;
wire n_552;
wire n_554;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_526;
wire n_485;
wire n_4038;
wire n_272;
wire n_271;
wire n_4043;
wire n_287;
wire n_286;
wire n_4047;
wire n_4048;
wire n_432;
wire n_431;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_550;
wire n_532;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_531;
wire n_4084;
wire n_4085;
wire n_484;
wire n_4087;
wire n_440;
wire n_427;
wire n_4092;
wire n_277;
wire n_270;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_331;
wire n_319;
wire n_4122;
wire n_375;
wire n_359;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4405;
wire n_4392;
wire n_4166;
wire n_4181;
wire n_4182;
wire n_415;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_315;
wire n_260;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_426;
wire n_416;
wire n_421;
wire n_417;
wire n_4213;
wire n_4473;
wire n_4470;
wire n_4219;
wire n_225;
wire n_224;
wire n_4223;
wire n_4435;
wire n_4434;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4452;
wire n_4247;
wire n_4449;
wire n_4249;
wire n_4451;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4384;
wire n_4382;
wire n_4262;
wire n_316;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4457;
wire n_4448;
wire n_4283;
wire n_4439;
wire n_4444;
wire n_4443;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4431;
wire n_4437;
wire n_4317;
wire n_4318;
wire n_4380;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_205;
wire n_204;
wire n_4336;
wire n_4339;
wire n_4516;
wire n_4340;
wire n_4341;
wire n_222;
wire n_4343;
wire n_176;
wire n_170;
wire n_4348;
wire n_196;
wire n_195;
wire n_4352;
wire n_4355;
wire n_4512;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4419;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4513;
wire n_4511;
wire n_4383;
wire n_190;
wire n_169;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_221;
wire n_4397;
wire n_4398;
wire n_4438;
wire n_4399;
wire n_4447;
wire n_4420;
wire n_4430;
wire n_4400;
wire n_4401;
wire n_151;
wire n_150;
wire n_4407;
wire n_142;
wire n_141;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_157;
wire n_156;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4496;
wire n_4491;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_130;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4483;
wire n_4482;
wire n_4479;
wire n_4549;
wire n_4551;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4565;
wire n_4571;
wire n_4521;
wire n_4481;
wire n_4524;
wire n_4532;
wire n_4552;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4575;
wire n_4616;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_110;
wire n_109;
wire n_4570;
wire n_102;
wire n_101;
wire n_4576;
wire n_106;
wire n_4577;
wire n_4601;
wire n_4613;
wire n_4600;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4593;
wire n_4581;
wire n_4595;
wire n_4582;
wire n_4596;
wire n_4594;
wire n_4583;
wire n_4584;
wire n_4597;
wire n_4615;
wire n_4599;
wire n_4614;
wire n_4585;
wire n_4586;
wire n_4617;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_107;
wire n_96;
wire n_4598;
wire n_87;
wire n_86;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_81;
wire n_85;
wire n_4624;
wire n_92;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_80;
wire n_4629;
wire n_79;
wire n_4631;
wire n_0;
wire n_1;
wire n_4618;
wire n_2;
wire n_4;
wire n_5;
wire n_4620;
wire n_129;
wire n_125;
wire n_6;
wire n_91;
wire n_7;
wire n_8;
wire n_52;
wire n_59;
wire n_62;
wire n_54;
wire n_53;
wire n_57;
wire n_56;
wire n_58;
wire n_60;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_83;
wire n_82;
wire n_123;
wire n_84;
wire n_128;
wire n_89;
wire n_122;
wire n_88;
wire n_105;
wire n_124;
wire n_100;
wire n_99;
wire n_97;
wire n_98;
wire n_104;
wire n_103;
wire n_111;
wire n_113;
wire n_112;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_126;
wire n_114;
wire n_168;
wire n_131;
wire n_132;
wire n_136;
wire n_135;
wire n_133;
wire n_138;
wire n_137;
wire n_146;
wire n_140;
wire n_145;
wire n_139;
wire n_144;
wire n_143;
wire n_203;
wire n_147;
wire n_149;
wire n_148;
wire n_155;
wire n_154;
wire n_167;
wire n_165;
wire n_152;
wire n_153;
wire n_158;
wire n_164;
wire n_191;
wire n_178;
wire n_177;
wire n_174;
wire n_172;
wire n_171;
wire n_173;
wire n_175;
wire n_188;
wire n_187;
wire n_186;
wire n_185;
wire n_182;
wire n_180;
wire n_179;
wire n_181;
wire n_184;
wire n_183;
wire n_219;
wire n_214;
wire n_189;
wire n_193;
wire n_192;
wire n_202;
wire n_201;
wire n_194;
wire n_208;
wire n_206;
wire n_200;
wire n_207;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_230;
wire n_228;
wire n_223;
wire n_226;
wire n_227;
wire n_238;
wire n_237;
wire n_254;
wire n_246;
wire n_239;
wire n_258;
wire n_256;
wire n_255;
wire n_257;
wire n_302;
wire n_261;
wire n_269;
wire n_262;
wire n_266;
wire n_264;
wire n_263;
wire n_265;
wire n_268;
wire n_267;
wire n_279;
wire n_278;
wire n_276;
wire n_275;
wire n_273;
wire n_274;
wire n_301;
wire n_300;
wire n_280;
wire n_284;
wire n_283;
wire n_310;
wire n_285;
wire n_305;
wire n_303;
wire n_304;
wire n_308;
wire n_307;
wire n_313;
wire n_312;
wire n_311;
wire n_309;
wire n_318;
wire n_317;
wire n_333;
wire n_381;
wire n_376;
wire n_328;
wire n_327;
wire n_330;
wire n_329;
wire n_338;
wire n_334;
wire n_340;
wire n_339;
wire n_358;
wire n_360;
wire n_363;
wire n_361;
wire n_372;
wire n_362;
wire n_373;
wire n_392;
wire n_390;
wire n_382;
wire n_384;
wire n_383;
wire n_385;
wire n_388;
wire n_394;
wire n_393;
wire n_399;
wire n_398;
wire n_395;
wire n_397;
wire n_418;
wire n_420;
wire n_419;
wire n_481;
wire n_423;
wire n_422;
wire n_483;
wire n_425;
wire n_424;
wire n_460;
wire n_430;
wire n_428;
wire n_429;
wire n_439;
wire n_438;
wire n_437;
wire n_436;
wire n_480;
wire n_433;
wire n_452;
wire n_450;
wire n_449;
wire n_448;
wire n_441;
wire n_447;
wire n_446;
wire n_444;
wire n_479;
wire n_451;
wire n_459;
wire n_457;
wire n_456;
wire n_458;
wire n_528;
wire n_527;
wire n_487;
wire n_489;
wire n_488;
wire n_518;
wire n_525;
wire n_496;
wire n_494;
wire n_499;
wire n_497;
wire n_498;
wire n_508;
wire n_507;
wire n_516;
wire n_517;
wire n_523;
wire n_524;
wire n_533;
wire n_543;
wire n_534;
wire n_547;
wire n_545;
wire n_549;
wire n_548;
wire n_560;
wire n_558;
wire n_557;
wire n_563;
wire n_562;
wire n_573;
wire n_572;
wire n_564;
wire n_569;
wire n_568;
wire n_586;
wire n_587;
wire n_576;
wire n_581;
wire n_582;
wire n_592;
wire n_591;
wire n_600;
wire n_593;
wire n_639;
wire n_632;
wire n_599;
wire n_598;
wire n_595;
wire n_594;
wire n_596;
wire n_597;
wire n_608;
wire n_601;
wire n_605;
wire n_603;
wire n_602;
wire n_667;
wire n_604;
wire n_607;
wire n_606;
wire n_629;
wire n_627;
wire n_609;
wire n_610;
wire n_628;
wire n_631;
wire n_630;
wire n_637;
wire n_635;
wire n_633;
wire n_634;
wire n_636;
wire n_638;
wire n_669;
wire n_641;
wire n_640;
wire n_644;
wire n_643;
wire n_642;
wire n_646;
wire n_645;
wire n_668;
wire n_647;
wire n_656;
wire n_649;
wire n_653;
wire n_651;
wire n_650;
wire n_652;
wire n_655;
wire n_654;
wire n_661;
wire n_657;
wire n_671;
wire n_658;
wire n_670;
wire n_660;
wire n_659;
wire n_665;
wire n_663;
wire n_662;
wire n_664;
wire n_666;
wire n_672;
wire n_673;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_704;
wire n_705;
wire n_706;
wire n_708;
wire n_712;
wire n_716;
wire n_854;
wire n_855;
wire n_748;
wire n_747;
wire n_722;
wire n_723;
wire n_738;
wire n_731;
wire n_726;
wire n_727;
wire n_773;
wire n_849;
wire n_728;
wire n_730;
wire n_729;
wire n_740;
wire n_739;
wire n_743;
wire n_805;
wire n_741;
wire n_787;
wire n_745;
wire n_742;
wire n_796;
wire n_744;
wire n_746;
wire n_750;
wire n_749;
wire n_752;
wire n_751;
wire n_857;
wire n_755;
wire n_753;
wire n_754;
wire n_878;
wire n_760;
wire n_759;
wire n_768;
wire n_758;
wire n_762;
wire n_761;
wire n_765;
wire n_764;
wire n_882;
wire n_859;
wire n_766;
wire n_809;
wire n_807;
wire n_806;
wire n_769;
wire n_795;
wire n_794;
wire n_793;
wire n_770;
wire n_785;
wire n_784;
wire n_786;
wire n_792;
wire n_800;
wire n_797;
wire n_804;
wire n_802;
wire n_801;
wire n_798;
wire n_799;
wire n_803;
wire n_879;
wire n_808;
wire n_822;
wire n_821;
wire n_810;
wire n_844;
wire n_843;
wire n_842;
wire n_834;
wire n_815;
wire n_814;
wire n_813;
wire n_811;
wire n_812;
wire n_816;
wire n_824;
wire n_823;
wire n_828;
wire n_827;
wire n_826;
wire n_825;
wire n_829;
wire n_832;
wire n_858;
wire n_830;
wire n_831;
wire n_835;
wire n_841;
wire n_837;
wire n_836;
wire n_839;
wire n_838;
wire n_848;
wire n_847;
wire n_845;
wire n_851;
wire n_865;
wire n_850;
wire n_846;
wire n_880;
wire n_852;
wire n_1585;
wire n_941;
wire n_890;
wire n_889;
wire n_887;
wire n_885;
wire n_888;
wire n_886;
wire n_900;
wire n_891;
wire n_937;
wire n_936;
wire n_903;
wire n_896;
wire n_1095;
wire n_894;
wire n_898;
wire n_897;
wire n_1100;
wire n_1099;
wire n_1085;
wire n_1084;
wire n_902;
wire n_901;
wire n_1052;
wire n_1051;
wire n_904;
wire n_920;
wire n_919;
wire n_918;
wire n_905;
wire n_913;
wire n_912;
wire n_911;
wire n_906;
wire n_907;
wire n_910;
wire n_909;
wire n_908;
wire n_1451;
wire n_915;
wire n_914;
wire n_1123;
wire n_917;
wire n_916;
wire n_925;
wire n_924;
wire n_922;
wire n_921;
wire n_923;
wire n_1579;
wire n_1577;
wire n_1576;
wire n_935;
wire n_929;
wire n_1582;
wire n_1580;
wire n_1250;
wire n_1246;
wire n_1245;
wire n_939;
wire n_938;
wire n_1109;
wire n_1103;
wire n_1082;
wire n_1081;
wire n_1018;
wire n_948;
wire n_946;
wire n_944;
wire n_1025;
wire n_950;
wire n_949;
wire n_1009;
wire n_1015;
wire n_1010;
wire n_1000;
wire n_1002;
wire n_1001;
wire n_957;
wire n_954;
wire n_953;
wire n_1044;
wire n_997;
wire n_983;
wire n_1022;
wire n_989;
wire n_1036;
wire n_1035;
wire n_1004;
wire n_1131;
wire n_1003;
wire n_1127;
wire n_1008;
wire n_1007;
wire n_1012;
wire n_1011;
wire n_1023;
wire n_1028;
wire n_1026;
wire n_1027;
wire n_1037;
wire n_1124;
wire n_1043;
wire n_1047;
wire n_1045;
wire n_1046;
wire n_1102;
wire n_1080;
wire n_1079;
wire n_1050;
wire n_1054;
wire n_1053;
wire n_1058;
wire n_1057;
wire n_1055;
wire n_1076;
wire n_1061;
wire n_1060;
wire n_1126;
wire n_1078;
wire n_1056;
wire n_1059;
wire n_1075;
wire n_1077;
wire n_1097;
wire n_1093;
wire n_1098;
wire n_1094;
wire n_1083;
wire n_1086;
wire n_1096;
wire n_1101;
wire n_1122;
wire n_1112;
wire n_1132;
wire n_1217;
wire n_1216;
wire n_1215;
wire n_1138;
wire n_1141;
wire n_1140;
wire n_1151;
wire n_1145;
wire n_1144;
wire n_1150;
wire n_1149;
wire n_1166;
wire n_1165;
wire n_1157;
wire n_1168;
wire n_1167;
wire n_1182;
wire n_1181;
wire n_1183;
wire n_1169;
wire n_1201;
wire n_1200;
wire n_1187;
wire n_1179;
wire n_1180;
wire n_1186;
wire n_1185;
wire n_1184;
wire n_1190;
wire n_1189;
wire n_1188;
wire n_1198;
wire n_1199;
wire n_1203;
wire n_1202;
wire n_1208;
wire n_1206;
wire n_1205;
wire n_1204;
wire n_1213;
wire n_1211;
wire n_1210;
wire n_1207;
wire n_1209;
wire n_1212;
wire n_1214;
wire n_1224;
wire n_1223;
wire n_1313;
wire n_1228;
wire n_1227;
wire n_1280;
wire n_1226;
wire n_1243;
wire n_1241;
wire n_1240;
wire n_1229;
wire n_1232;
wire n_1231;
wire n_1230;
wire n_1239;
wire n_1238;
wire n_1252;
wire n_1251;
wire n_1244;
wire n_1247;
wire n_1542;
wire n_1254;
wire n_1253;
wire n_1284;
wire n_1283;
wire n_1282;
wire n_1281;
wire n_1295;
wire n_1296;
wire n_1285;
wire n_1290;
wire n_1289;
wire n_1286;
wire n_1348;
wire n_1288;
wire n_1287;
wire n_1292;
wire n_1291;
wire n_3272;
wire n_3270;
wire n_3269;
wire n_1293;
wire n_3255;
wire n_3254;
wire n_3107;
wire n_1432;
wire n_1298;
wire n_1297;
wire n_1294;
wire n_1305;
wire n_1304;
wire n_1300;
wire n_1311;
wire n_1310;
wire n_1309;
wire n_1308;
wire n_1303;
wire n_1302;
wire n_1301;
wire n_3097;
wire n_1307;
wire n_1306;
wire n_3250;
wire n_3284;
wire n_3281;
wire n_3280;
wire n_3279;
wire n_3277;
wire n_1315;
wire n_1314;
wire n_1343;
wire n_1342;
wire n_1341;
wire n_1316;
wire n_1326;
wire n_1325;
wire n_1324;
wire n_1317;
wire n_1331;
wire n_1330;
wire n_1332;
wire n_1327;
wire n_1340;
wire n_1339;
wire n_1334;
wire n_1333;
wire n_1347;
wire n_1346;
wire n_1345;
wire n_1344;
wire n_1356;
wire n_1360;
wire n_1358;
wire n_1393;
wire n_1392;
wire n_1419;
wire n_1391;
wire n_1410;
wire n_1409;
wire n_1394;
wire n_1398;
wire n_1396;
wire n_1395;
wire n_1400;
wire n_1399;
wire n_1408;
wire n_1412;
wire n_1411;
wire n_1418;
wire n_1417;
wire n_1416;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1547;
wire n_1422;
wire n_1421;
wire n_1420;
wire n_1424;
wire n_1423;
wire n_1445;
wire n_1443;
wire n_1442;
wire n_1425;
wire n_1435;
wire n_1434;
wire n_1433;
wire n_1426;
wire n_1427;
wire n_1431;
wire n_1429;
wire n_1428;
wire n_1430;
wire n_1436;
wire n_1440;
wire n_1439;
wire n_1441;
wire n_1537;
wire n_1536;
wire n_1535;
wire n_1488;
wire n_1446;
wire n_1463;
wire n_1462;
wire n_1447;
wire n_1456;
wire n_1452;
wire n_1450;
wire n_1453;
wire n_1460;
wire n_1465;
wire n_1464;
wire n_1470;
wire n_1467;
wire n_1466;
wire n_1482;
wire n_1474;
wire n_1472;
wire n_1480;
wire n_1473;
wire n_1487;
wire n_1511;
wire n_1489;
wire n_1512;
wire n_1513;
wire n_1546;
wire n_1545;
wire n_1544;
wire n_1543;
wire n_1538;
wire n_1540;
wire n_1650;
wire n_1560;
wire n_1562;
wire n_1561;
wire n_1564;
wire n_1648;
wire n_1563;
wire n_1567;
wire n_1565;
wire n_1566;
wire n_1570;
wire n_1569;
wire n_1568;
wire n_1575;
wire n_1574;
wire n_1586;
wire n_1573;
wire n_1572;
wire n_1571;
wire n_1581;
wire n_1593;
wire n_1592;
wire n_1606;
wire n_1591;
wire n_1598;
wire n_1595;
wire n_1594;
wire n_1600;
wire n_1599;
wire n_1597;
wire n_1646;
wire n_1603;
wire n_1641;
wire n_1640;
wire n_1639;
wire n_1607;
wire n_1635;
wire n_1634;
wire n_1633;
wire n_1637;
wire n_1636;
wire n_1638;
wire n_1647;
wire n_1645;
wire n_1644;
wire n_1643;
wire n_3391;
wire n_1642;
wire n_1652;
wire n_1651;
wire n_1717;
wire n_1716;
wire n_1662;
wire n_1677;
wire n_1663;
wire n_1664;
wire n_1692;
wire n_1689;
wire n_1678;
wire n_1710;
wire n_1709;
wire n_1708;
wire n_1707;
wire n_1684;
wire n_1681;
wire n_1680;
wire n_1679;
wire n_1682;
wire n_1685;
wire n_1694;
wire n_1693;
wire n_1699;
wire n_1698;
wire n_1697;
wire n_1706;
wire n_1705;
wire n_1704;
wire n_1703;
wire n_1701;
wire n_1700;
wire n_1702;
wire n_1720;
wire n_1722;
wire n_1721;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1798;
wire n_1800;
wire n_1799;
wire n_1802;
wire n_1866;
wire n_1865;
wire n_1864;
wire n_1856;
wire n_1804;
wire n_1803;
wire n_1805;
wire n_1808;
wire n_1825;
wire n_1807;
wire n_1810;
wire n_1809;
wire n_1819;
wire n_1813;
wire n_1812;
wire n_1811;
wire n_1824;
wire n_1823;
wire n_1821;
wire n_1820;
wire n_1822;
wire n_1835;
wire n_1834;
wire n_1827;
wire n_1826;
wire n_1833;
wire n_1831;
wire n_1828;
wire n_1832;
wire n_1829;
wire n_1837;
wire n_1836;
wire n_1842;
wire n_1840;
wire n_1839;
wire n_1838;
wire n_1894;
wire n_1845;
wire n_1844;
wire n_1841;
wire n_1843;
wire n_1847;
wire n_1846;
wire n_1857;
wire n_1858;
wire n_1862;
wire n_1861;
wire n_1860;
wire n_1859;
wire n_1863;
wire n_1868;
wire n_1867;
wire n_1889;
wire n_1869;
wire n_1888;
wire n_1887;
wire n_1886;
wire n_1870;
wire n_1893;
wire n_1892;
wire n_1891;
wire n_1890;
wire n_1895;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1904;
wire n_1905;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1939;
wire n_1933;
wire n_1935;
wire n_1934;
wire n_1937;
wire n_1936;
wire n_1938;
wire n_1960;
wire n_1940;
wire n_1945;
wire n_1944;
wire n_1947;
wire n_1946;
wire n_1948;
wire n_1961;
wire n_1963;
wire n_1962;
wire n_1964;
wire n_1994;
wire n_1966;
wire n_1972;
wire n_1967;
wire n_1970;
wire n_1968;
wire n_1969;
wire n_2013;
wire n_1971;
wire n_1974;
wire n_1973;
wire n_2010;
wire n_2008;
wire n_1985;
wire n_1984;
wire n_1975;
wire n_1982;
wire n_1981;
wire n_1993;
wire n_1986;
wire n_1990;
wire n_1989;
wire n_2003;
wire n_1995;
wire n_2002;
wire n_2001;
wire n_2011;
wire n_2007;
wire n_2005;
wire n_2036;
wire n_2009;
wire n_2035;
wire n_2015;
wire n_2014;
wire n_2012;
wire n_2016;
wire n_2090;
wire n_2048;
wire n_2047;
wire n_2040;
wire n_2043;
wire n_2042;
wire n_2041;
wire n_2074;
wire n_2073;
wire n_2045;
wire n_2044;
wire n_2069;
wire n_2068;
wire n_2101;
wire n_2046;
wire n_2102;
wire n_2100;
wire n_2050;
wire n_2049;
wire n_2053;
wire n_2052;
wire n_2051;
wire n_2066;
wire n_2060;
wire n_2055;
wire n_2054;
wire n_2061;
wire n_2063;
wire n_2062;
wire n_2094;
wire n_2098;
wire n_2097;
wire n_2072;
wire n_2067;
wire n_2065;
wire n_2064;
wire n_2071;
wire n_2070;
wire n_2117;
wire n_2076;
wire n_2075;
wire n_2081;
wire n_2080;
wire n_2079;
wire n_2092;
wire n_2091;
wire n_2106;
wire n_2105;
wire n_2093;
wire n_2096;
wire n_2095;
wire n_2099;
wire n_2103;
wire n_2104;
wire n_2118;
wire n_2116;
wire n_2115;
wire n_2108;
wire n_2107;
wire n_2146;
wire n_2141;
wire n_2109;
wire n_2168;
wire n_2111;
wire n_2114;
wire n_2112;
wire n_2113;
wire n_2129;
wire n_2127;
wire n_2126;
wire n_2120;
wire n_2125;
wire n_2124;
wire n_2128;
wire n_2133;
wire n_2138;
wire n_2132;
wire n_2135;
wire n_2134;
wire n_2139;
wire n_2148;
wire n_2147;
wire n_2149;
wire n_2167;
wire n_2166;
wire n_2165;
wire n_2161;
wire n_2163;
wire n_2162;
wire n_2164;
wire n_2169;
wire n_2173;
wire n_2172;
wire n_2179;
wire n_2176;
wire n_2175;
wire n_2178;
wire n_2181;
wire n_2180;
wire n_2185;
wire n_2184;
wire n_2183;
wire n_2191;
wire n_2192;
wire n_2189;
wire n_2193;
wire n_2190;
wire n_2194;
wire n_2197;
wire n_2201;
wire n_2199;
wire n_2198;
wire n_2200;
wire n_2202;
wire n_2234;
wire n_2224;
wire n_2215;
wire n_2222;
wire n_2216;
wire n_2220;
wire n_2218;
wire n_2217;
wire n_2219;
wire n_2245;
wire n_2221;
wire n_2223;
wire n_2226;
wire n_2225;
wire n_2230;
wire n_2228;
wire n_2227;
wire n_2229;
wire n_2232;
wire n_2231;
wire n_2236;
wire n_2235;
wire n_2242;
wire n_2238;
wire n_2237;
wire n_2243;
wire n_2239;
wire n_2240;
wire n_2244;
wire n_2251;
wire n_2250;
wire n_2253;
wire n_2255;
wire n_2252;
wire n_2254;
wire n_2257;
wire n_2258;
wire n_2264;
wire n_2263;
wire n_2262;
wire n_2261;
wire n_2276;
wire n_2275;
wire n_2265;
wire n_2318;
wire n_2267;
wire n_2268;
wire n_2266;
wire n_2269;
wire n_2273;
wire n_2271;
wire n_2270;
wire n_2272;
wire n_2285;
wire n_2274;
wire n_2278;
wire n_2277;
wire n_2284;
wire n_2283;
wire n_2280;
wire n_2279;
wire n_2281;
wire n_2282;
wire n_2315;
wire n_2313;
wire n_2317;
wire n_2316;
wire n_2322;
wire n_2324;
wire n_2323;
wire n_2343;
wire n_2339;
wire n_2326;
wire n_2348;
wire n_2347;
wire n_2346;
wire n_2330;
wire n_2341;
wire n_2340;
wire n_2342;
wire n_2345;
wire n_2344;
wire n_2352;
wire n_2351;
wire n_2354;
wire n_2353;
wire n_2360;
wire n_2406;
wire n_2358;
wire n_2369;
wire n_2361;
wire n_2409;
wire n_2403;
wire n_2402;
wire n_2370;
wire n_2368;
wire n_2382;
wire n_2376;
wire n_2378;
wire n_2377;
wire n_2395;
wire n_2400;
wire n_2399;
wire n_2392;
wire n_2385;
wire n_2384;
wire n_2383;
wire n_2393;
wire n_2398;
wire n_2394;
wire n_2396;
wire n_2397;
wire n_2407;
wire n_2404;
wire n_2408;
wire n_2405;
wire n_2401;
wire n_2479;
wire n_2455;
wire n_2454;
wire n_2417;
wire n_2416;
wire n_2464;
wire n_2463;
wire n_2425;
wire n_2469;
wire n_2468;
wire n_2419;
wire n_2427;
wire n_2426;
wire n_2500;
wire n_2431;
wire n_2428;
wire n_2438;
wire n_2437;
wire n_2435;
wire n_2452;
wire n_2440;
wire n_2462;
wire n_2461;
wire n_2460;
wire n_2467;
wire n_2466;
wire n_2465;
wire n_2523;
wire n_2518;
wire n_2513;
wire n_2509;
wire n_2472;
wire n_2470;
wire n_2473;
wire n_2471;
wire n_2499;
wire n_2497;
wire n_2496;
wire n_2504;
wire n_2492;
wire n_2481;
wire n_2480;
wire n_2525;
wire n_2526;
wire n_2485;
wire n_2487;
wire n_2486;
wire n_2495;
wire n_2491;
wire n_2488;
wire n_2507;
wire n_2493;
wire n_2494;
wire n_2498;
wire n_2503;
wire n_2505;
wire n_2517;
wire n_2508;
wire n_2511;
wire n_2510;
wire n_2512;
wire n_2520;
wire n_2519;
wire n_2522;
wire n_2521;
wire n_2528;
wire n_2527;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2553;
wire n_2554;
wire n_2556;
wire n_2561;
wire n_2573;
wire n_2579;
wire n_2580;
wire n_2589;
wire n_2588;
wire n_2608;
wire n_2586;
wire n_2610;
wire n_2611;
wire n_2598;
wire n_2597;
wire n_2590;
wire n_2600;
wire n_2599;
wire n_2601;
wire n_2605;
wire n_2620;
wire n_2617;
wire n_2609;
wire n_2625;
wire n_2628;
wire n_2624;
wire n_2623;
wire n_2616;
wire n_2618;
wire n_2619;
wire n_2621;
wire n_2627;
wire n_2626;
wire n_2632;
wire n_2634;
wire n_2653;
wire n_2645;
wire n_2649;
wire n_2646;
wire n_2648;
wire n_2652;
wire n_2655;
wire n_2665;
wire n_2658;
wire n_2664;
wire n_2660;
wire n_2659;
wire n_2661;
wire n_2662;
wire n_2670;
wire n_2666;
wire n_2669;
wire n_2668;
wire n_2667;
wire n_2674;
wire n_2673;
wire n_2672;
wire n_2671;
wire n_2678;
wire n_2677;
wire n_2693;
wire n_2684;
wire n_2683;
wire n_2687;
wire n_2686;
wire n_2689;
wire n_2691;
wire n_2690;
wire n_2688;
wire n_2695;
wire n_2694;
wire n_2696;
wire n_2703;
wire n_2701;
wire n_2702;
wire n_2705;
wire n_2704;
wire n_2709;
wire n_2707;
wire n_2708;
wire n_2711;
wire n_2710;
wire n_2713;
wire n_2743;
wire n_2742;
wire n_2716;
wire n_2718;
wire n_2738;
wire n_2739;
wire n_2753;
wire n_2752;
wire n_2744;
wire n_2748;
wire n_2747;
wire n_2749;
wire n_2757;
wire n_2756;
wire n_2773;
wire n_2772;
wire n_2762;
wire n_2758;
wire n_2761;
wire n_2763;
wire n_2770;
wire n_2767;
wire n_2766;
wire n_2768;
wire n_2769;
wire n_2782;
wire n_2776;
wire n_2774;
wire n_2783;
wire n_2787;
wire n_2777;
wire n_2775;
wire n_2788;
wire n_2784;
wire n_2786;
wire n_2785;
wire n_2805;
wire n_2795;
wire n_2836;
wire n_2835;
wire n_2797;
wire n_2796;
wire n_2847;
wire n_2846;
wire n_2841;
wire n_2848;
wire n_2842;
wire n_2801;
wire n_2812;
wire n_2811;
wire n_2803;
wire n_2802;
wire n_2821;
wire n_2817;
wire n_2816;
wire n_2904;
wire n_2909;
wire n_2908;
wire n_2810;
wire n_2813;
wire n_2891;
wire n_2818;
wire n_2820;
wire n_2824;
wire n_2822;
wire n_2823;
wire n_2833;
wire n_2829;
wire n_2828;
wire n_2830;
wire n_2838;
wire n_2834;
wire n_2837;
wire n_2839;
wire n_2845;
wire n_2840;
wire n_2844;
wire n_2843;
wire n_2849;
wire n_2874;
wire n_2876;
wire n_2875;
wire n_2896;
wire n_2895;
wire n_2877;
wire n_2883;
wire n_2882;
wire n_2889;
wire n_2898;
wire n_2901;
wire n_2911;
wire n_2907;
wire n_2910;
wire n_2936;
wire n_2928;
wire n_2930;
wire n_2929;
wire n_2932;
wire n_2931;
wire n_2998;
wire n_2935;
wire n_2960;
wire n_2937;
wire n_2946;
wire n_2945;
wire n_2938;
wire n_2943;
wire n_2939;
wire n_2942;
wire n_2944;
wire n_2948;
wire n_2947;
wire n_2958;
wire n_2953;
wire n_2951;
wire n_2952;
wire n_2956;
wire n_2957;
wire n_2975;
wire n_2976;
wire n_2962;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2969;
wire n_2971;
wire n_2977;
wire n_2990;
wire n_2980;
wire n_3011;
wire n_3009;
wire n_3013;
wire n_3012;
wire n_3019;
wire n_3018;
wire n_3031;
wire n_3017;
wire n_3024;
wire n_3022;
wire n_3020;
wire n_3030;
wire n_3026;
wire n_3025;
wire n_3023;
wire n_3029;
wire n_3039;
wire n_3038;
wire n_3033;
wire n_3032;
wire n_3051;
wire n_3043;
wire n_3042;
wire n_3049;
wire n_3050;
wire n_3098;
wire n_3073;
wire n_3096;
wire n_3095;
wire n_3075;
wire n_3074;
wire n_3150;
wire n_3101;
wire n_3149;
wire n_3099;
wire n_3131;
wire n_3102;
wire n_3106;
wire n_3104;
wire n_3103;
wire n_3105;
wire n_3144;
wire n_3132;
wire n_3136;
wire n_3133;
wire n_3137;
wire n_3134;
wire n_3148;
wire n_3147;
wire n_3146;
wire n_3145;
wire n_3156;
wire n_3151;
wire n_3155;
wire n_3153;
wire n_3152;
wire n_3154;
wire n_3174;
wire n_3157;
wire n_3172;
wire n_3170;
wire n_3171;
wire n_3169;
wire n_3178;
wire n_3177;
wire n_3176;
wire n_3175;
wire n_3198;
wire n_3196;
wire n_3184;
wire n_3183;
wire n_3194;
wire n_3193;
wire n_3201;
wire n_3205;
wire n_3204;
wire n_3207;
wire n_3209;
wire n_3208;
wire n_3217;
wire n_3213;
wire n_3216;
wire n_3232;
wire n_3237;
wire n_3245;
wire n_3244;
wire n_3285;
wire n_3238;
wire n_3249;
wire n_3248;
wire n_3274;
wire n_3251;
wire n_3252;
wire n_3271;
wire n_3276;
wire n_3275;
wire n_3278;
wire n_3283;
wire n_3287;
wire n_3286;
wire n_3292;
wire n_3288;
wire n_3290;
wire n_3289;
wire n_3293;
wire n_3326;
wire n_3325;
wire n_3324;
wire n_3296;
wire n_3299;
wire n_3298;
wire n_3303;
wire n_3302;
wire n_3314;
wire n_3313;
wire n_3319;
wire n_3318;
wire n_3431;
wire n_3347;
wire n_3346;
wire n_3350;
wire n_3352;
wire n_3351;
wire n_3358;
wire n_3357;
wire n_3356;
wire n_3354;
wire n_3355;
wire n_3432;
wire n_3372;
wire n_3371;
wire n_3360;
wire n_3359;
wire n_3394;
wire n_3393;
wire n_3392;
wire n_3382;
wire n_3451;
wire n_3433;
wire n_3370;
wire n_3361;
wire n_3374;
wire n_3373;
wire n_3378;
wire n_3387;
wire n_3386;
wire n_3383;
wire n_3390;
wire n_3399;
wire n_3398;
wire n_3397;
wire n_3412;
wire n_3411;
wire n_3410;
wire n_3409;
wire n_3430;
wire n_3429;
wire n_3428;
wire n_3413;
wire n_3414;
wire n_3424;
wire n_3423;
wire n_3415;
wire n_3416;
wire n_3420;
wire n_3422;
wire n_3421;
wire n_3426;
wire n_3425;
wire n_3452;
wire n_3456;
wire n_3458;
wire n_3457;
wire n_3460;
wire n_3462;
wire n_3461;
wire n_3466;
wire n_3465;
wire n_3470;
wire n_3472;
wire n_3471;
wire n_3487;
wire n_3486;
wire n_3474;
wire n_3479;
wire n_3478;
wire n_3476;
wire n_3482;
wire n_3481;
wire n_3484;
wire n_3483;
wire n_3516;
wire n_3508;
wire n_3498;
wire n_3497;
wire n_3493;
wire n_3492;
wire n_3506;
wire n_3501;
wire n_3512;
wire n_3511;
wire n_3525;
wire n_3519;
wire n_3542;
wire n_3541;
wire n_3539;
wire n_3544;
wire n_3545;
wire n_3563;
wire n_3570;
wire n_3569;
wire n_3586;
wire n_3590;
wire n_3589;
wire n_3587;
wire n_3585;
wire n_3584;
wire n_3603;
wire n_3601;
wire n_3598;
wire n_3591;
wire n_3595;
wire n_3593;
wire n_3592;
wire n_3594;
wire n_3597;
wire n_3612;
wire n_3611;
wire n_3609;
wire n_3608;
wire n_3607;
wire n_3606;
wire n_3621;
wire n_3619;
wire n_3613;
wire n_3623;
wire n_3620;
wire n_3618;
wire n_3622;
wire n_3625;
wire n_3722;
wire n_3630;
wire n_3629;
wire n_3641;
wire n_3638;
wire n_3637;
wire n_3632;
wire n_3631;
wire n_3777;
wire n_3675;
wire n_3640;
wire n_3639;
wire n_3636;
wire n_3679;
wire n_3678;
wire n_3669;
wire n_3674;
wire n_3673;
wire n_3676;
wire n_3718;
wire n_3717;
wire n_3682;
wire n_3683;
wire n_3687;
wire n_3697;
wire n_3724;
wire n_3723;
wire n_3736;
wire n_3725;
wire n_3735;
wire n_3734;
wire n_3731;
wire n_3733;
wire n_3782;
wire n_3737;
wire n_3776;
wire n_3745;
wire n_3739;
wire n_3775;
wire n_3787;
wire n_3785;
wire n_3783;
wire n_3784;
wire n_3786;
wire n_3797;
wire n_3940;
wire n_3939;
wire n_3941;
wire n_3938;
wire n_3822;
wire n_3817;
wire n_3803;
wire n_3802;
wire n_3816;
wire n_3820;
wire n_3852;
wire n_3823;
wire n_3858;
wire n_3854;
wire n_3853;
wire n_3862;
wire n_3860;
wire n_3859;
wire n_3855;
wire n_3856;
wire n_3861;
wire n_3892;
wire n_3895;
wire n_3894;
wire n_3908;
wire n_3906;
wire n_3937;
wire n_3909;
wire n_3947;
wire n_3946;
wire n_3967;
wire n_3966;
wire n_4036;
wire n_4041;
wire n_4040;
wire n_3962;
wire n_4007;
wire n_4006;
wire n_3964;
wire n_3963;
wire n_4031;
wire n_4030;
wire n_4027;
wire n_4024;
wire n_3977;
wire n_3969;
wire n_4009;
wire n_3993;
wire n_3973;
wire n_3972;
wire n_3986;
wire n_3978;
wire n_3982;
wire n_3981;
wire n_3984;
wire n_3983;
wire n_3985;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_4134;
wire n_3992;
wire n_4008;
wire n_4029;
wire n_4010;
wire n_4026;
wire n_4025;
wire n_4033;
wire n_4032;
wire n_4089;
wire n_4088;
wire n_4039;
wire n_4037;
wire n_4044;
wire n_4096;
wire n_4083;
wire n_4059;
wire n_4049;
wire n_4045;
wire n_4046;
wire n_4053;
wire n_4052;
wire n_4158;
wire n_4064;
wire n_4063;
wire n_4066;
wire n_4093;
wire n_4091;
wire n_4090;
wire n_4113;
wire n_4095;
wire n_4094;
wire n_4108;
wire n_4107;
wire n_4111;
wire n_4110;
wire n_4116;
wire n_4114;
wire n_4115;
wire n_4124;
wire n_4156;
wire n_4155;
wire n_4120;
wire n_4121;
wire n_4127;
wire n_4125;
wire n_4126;
wire n_4131;
wire n_4130;
wire n_4132;
wire n_4151;
wire n_4153;
wire n_4152;
wire n_4161;
wire n_4349;
wire n_4193;
wire n_4167;
wire n_4176;
wire n_4174;
wire n_4171;
wire n_4170;
wire n_4172;
wire n_4173;
wire n_4178;
wire n_4177;
wire n_4187;
wire n_4237;
wire n_4179;
wire n_4191;
wire n_4274;
wire n_4189;
wire n_4180;
wire n_4188;
wire n_4190;
wire n_4243;
wire n_4195;
wire n_4194;
wire n_4199;
wire n_4198;
wire n_4215;
wire n_4214;
wire n_4217;
wire n_4216;
wire n_4200;
wire n_4226;
wire n_4224;
wire n_4222;
wire n_4225;
wire n_4240;
wire n_4239;
wire n_4236;
wire n_4235;
wire n_4258;
wire n_4257;
wire n_4246;
wire n_4254;
wire n_4255;
wire n_4273;
wire n_4260;
wire n_4271;
wire n_4272;
wire n_4278;
wire n_4277;
wire n_4281;
wire n_4284;
wire n_4297;
wire n_4368;
wire n_4369;
wire n_4299;
wire n_4298;
wire n_4314;
wire n_4313;
wire n_4300;
wire n_4309;
wire n_4308;
wire n_4310;
wire n_4366;
wire n_4365;
wire n_4315;
wire n_4333;
wire n_4332;
wire n_4379;
wire n_4320;
wire n_4338;
wire n_4347;
wire n_4342;
wire n_4337;
wire n_4346;
wire n_4354;
wire n_4385;
wire n_4381;
wire n_4387;
wire n_4386;
wire n_4389;
wire n_4388;
wire n_4406;
wire n_4411;
wire n_4409;
wire n_4391;
wire n_4390;
wire n_4418;
wire n_4416;
wire n_4402;
wire n_4396;
wire n_4404;
wire n_4403;
wire n_4412;
wire n_4408;
wire n_4410;
wire n_4417;
wire n_4433;
wire n_4432;
wire n_4474;
wire n_4436;
wire n_4475;
wire n_4446;
wire n_4445;
wire n_4458;
wire n_4450;
wire n_4455;
wire n_4453;
wire n_4476;
wire n_4454;
wire n_4477;
wire n_4456;
wire n_4478;
wire n_4460;
wire n_4459;
wire n_4472;
wire n_4471;
wire n_4480;
wire n_4484;
wire n_4517;
wire n_4486;
wire n_4485;
wire n_4488;
wire n_4487;
wire n_4507;
wire n_4497;
wire n_4490;
wire n_4489;
wire n_4492;
wire n_4495;
wire n_4494;
wire n_4493;
wire n_4508;
wire n_4515;
wire n_4514;
wire n_4510;
wire n_4509;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4522;
wire n_4523;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4550;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4619;
wire n_4630;
wire n_4621;
wire n_4623;
wire n_4622;


AOI22_X1 i_4687 (.ZN (n_4630), .A1 (n_84), .A2 (n_91), .B1 (n_83), .B2 (n_82));
NAND2_X1 i_4686 (.ZN (n_4623), .A1 (inputA[30]), .A2 (inputB[31]));
NAND2_X1 i_4685 (.ZN (n_4622), .A1 (inputA[31]), .A2 (inputB[30]));
XNOR2_X1 i_4684 (.ZN (n_4621), .A (n_4623), .B (n_4622));
NOR2_X1 i_4683 (.ZN (n_4620), .A1 (n_4630), .A2 (n_4621));
AOI21_X1 i_4682 (.ZN (n_4619), .A (n_4620), .B1 (n_4630), .B2 (n_4621));
INV_X1 i_4681 (.ZN (n_4618), .A (n_4619));
OAI21_X1 i_4680 (.ZN (n_4617), .A (n_4574), .B1 (n_4575), .B2 (n_4616));
XNOR2_X1 i_4679 (.ZN (n_4616), .A (n_4597), .B (n_4615));
XOR2_X1 i_4678 (.Z (n_4615), .A (n_4614), .B (n_4599));
XOR2_X1 i_4677 (.Z (n_4614), .A (n_4601), .B (n_4613));
NOR2_X1 i_4676 (.ZN (n_4613), .A1 (n_215), .A2 (n_882));
XNOR2_X1 i_4675 (.ZN (n_4601), .A (n_4600), .B (n_106));
NAND2_X1 i_4674 (.ZN (n_4600), .A1 (inputB[31]), .A2 (inputA[26]));
XNOR2_X1 i_4673 (.ZN (n_4599), .A (n_114), .B (n_116));
XNOR2_X1 i_4670 (.ZN (n_4597), .A (n_4593), .B (n_4596));
XNOR2_X1 i_4669 (.ZN (n_4596), .A (n_4594), .B (n_4595));
AOI21_X1 i_4668 (.ZN (n_4595), .A (n_4566), .B1 (n_4568), .B2 (n_4569));
OAI33_X1 i_4667 (.ZN (n_4594), .A1 (n_4557), .A2 (n_214), .A3 (n_882), .B1 (n_128)
    , .B2 (n_215), .B3 (n_4555));
AOI22_X1 i_4665 (.ZN (n_4593), .A1 (n_4525), .A2 (n_4529), .B1 (n_4523), .B2 (n_4518));
OAI21_X1 i_4664 (.ZN (n_4575), .A (n_4574), .B1 (n_4572), .B2 (n_4573));
NAND2_X1 i_4663 (.ZN (n_4574), .A1 (n_4572), .A2 (n_4573));
OAI21_X1 i_4662 (.ZN (n_4573), .A (n_4564), .B1 (n_4565), .B2 (n_4571));
AOI22_X1 i_4661 (.ZN (n_4572), .A1 (n_4532), .A2 (n_4552), .B1 (n_4530), .B2 (n_4531));
XNOR2_X1 i_4660 (.ZN (n_4571), .A (n_4568), .B (n_4569));
NOR2_X1 i_4659 (.ZN (n_4569), .A1 (n_127), .A2 (n_122));
NOR2_X1 i_4658 (.ZN (n_4568), .A1 (n_4566), .A2 (n_4567));
AOI22_X1 i_4657 (.ZN (n_4567), .A1 (inputB[27]), .A2 (inputA[29]), .B1 (inputB[26]), .B2 (inputA[30]));
NOR2_X1 i_4656 (.ZN (n_4566), .A1 (n_4519), .A2 (n_114));
OAI21_X1 i_4655 (.ZN (n_4565), .A (n_4564), .B1 (n_4554), .B2 (n_4563));
NAND2_X1 i_4654 (.ZN (n_4564), .A1 (n_4554), .A2 (n_4563));
XOR2_X1 i_4653 (.Z (n_4563), .A (n_4557), .B (n_4562));
NAND2_X1 i_4652 (.ZN (n_4562), .A1 (inputB[30]), .A2 (inputA[26]));
XNOR2_X1 i_4651 (.ZN (n_4557), .A (n_4555), .B (n_4556));
NAND2_X1 i_4650 (.ZN (n_4556), .A1 (inputB[29]), .A2 (inputA[27]));
NOR2_X1 i_4647 (.ZN (n_4555), .A1 (n_129), .A2 (n_483));
NAND2_X1 i_4645 (.ZN (n_4554), .A1 (n_4553), .A2 (n_4543));
INV_X1 i_4644 (.ZN (n_4553), .A (n_4547));
AOI22_X1 i_4643 (.ZN (n_4552), .A1 (n_4549), .A2 (n_4551), .B1 (n_4540), .B2 (n_4548));
XOR2_X1 i_4642 (.Z (n_4551), .A (n_4522), .B (n_4550));
NAND2_X1 i_4641 (.ZN (n_4550), .A1 (inputB[28]), .A2 (inputA[27]));
XOR2_X1 i_4640 (.Z (n_4549), .A (n_4540), .B (n_4548));
AOI21_X1 i_4639 (.ZN (n_4548), .A (n_4547), .B1 (n_4546), .B2 (n_4544));
NOR2_X1 i_4638 (.ZN (n_4547), .A1 (n_4544), .A2 (n_4546));
AOI22_X1 i_4637 (.ZN (n_4546), .A1 (n_4545), .A2 (n_4508), .B1 (n_4510), .B2 (n_4509));
INV_X1 i_4636 (.ZN (n_4545), .A (n_154));
OAI21_X1 i_4635 (.ZN (n_4544), .A (n_4543), .B1 (n_4542), .B2 (n_4541));
NAND2_X1 i_4634 (.ZN (n_4543), .A1 (n_4541), .A2 (n_4542));
NOR2_X1 i_4633 (.ZN (n_4542), .A1 (n_219), .A2 (n_124));
NAND2_X1 i_4632 (.ZN (n_4541), .A1 (inputB[24]), .A2 (inputA[31]));
XOR2_X1 i_4631 (.Z (n_4540), .A (n_4528), .B (n_4539));
NAND2_X1 i_4630 (.ZN (n_4539), .A1 (inputA[25]), .A2 (inputB[30]));
XOR2_X1 i_4629 (.Z (n_4532), .A (n_4530), .B (n_4531));
AOI22_X1 i_4628 (.ZN (n_4531), .A1 (n_4487), .A2 (n_4488), .B1 (n_4490), .B2 (n_4489));
XNOR2_X1 i_4627 (.ZN (n_4530), .A (n_4525), .B (n_4529));
OAI33_X1 i_4626 (.ZN (n_4529), .A1 (n_4528), .A2 (n_483), .A3 (n_882), .B1 (n_214)
    , .B2 (n_128), .B3 (n_4526));
XNOR2_X1 i_4625 (.ZN (n_4528), .A (n_4526), .B (n_4527));
NAND2_X1 i_4624 (.ZN (n_4527), .A1 (inputB[29]), .A2 (inputA[26]));
NOR2_X1 i_4623 (.ZN (n_4526), .A1 (n_585), .A2 (n_129));
XOR2_X1 i_4622 (.Z (n_4525), .A (n_4518), .B (n_4523));
OAI33_X1 i_4621 (.ZN (n_4523), .A1 (n_4522), .A2 (n_127), .A3 (n_215), .B1 (n_4495)
    , .B2 (n_126), .B3 (n_123));
XNOR2_X1 i_4620 (.ZN (n_4522), .A (n_4519), .B (n_4520));
NAND2_X1 i_4619 (.ZN (n_4520), .A1 (inputA[28]), .A2 (inputB[27]));
NAND2_X1 i_4617 (.ZN (n_4519), .A1 (inputA[29]), .A2 (inputB[26]));
NAND2_X1 i_4616 (.ZN (n_4518), .A1 (inputB[25]), .A2 (inputA[31]));
INV_X1 i_4615 (.ZN (n_4517), .A (n_168));
XNOR2_X1 i_4614 (.ZN (n_4516), .A (n_189), .B (n_155));
NAND2_X1 i_4613 (.ZN (n_4515), .A1 (inputB[22]), .A2 (inputA[31]));
OAI33_X1 i_4612 (.ZN (n_4514), .A1 (n_219), .A2 (n_215), .A3 (n_4516), .B1 (n_155)
    , .B2 (n_461), .B3 (n_122));
XOR2_X1 i_4611 (.Z (n_4513), .A (n_4515), .B (n_4514));
XNOR2_X1 i_4610 (.ZN (n_4512), .A (n_183), .B (n_167));
OAI33_X1 i_4609 (.ZN (n_4511), .A1 (n_585), .A2 (n_127), .A3 (n_4512), .B1 (n_167)
    , .B2 (n_483), .B3 (n_126));
NOR2_X1 i_4608 (.ZN (n_4510), .A1 (n_219), .A2 (n_123));
NAND2_X1 i_4607 (.ZN (n_4509), .A1 (inputB[23]), .A2 (inputA[31]));
XOR2_X1 i_4606 (.Z (n_4508), .A (n_4510), .B (n_4509));
AOI22_X1 i_4605 (.ZN (n_4507), .A1 (n_4515), .A2 (n_4514), .B1 (n_4513), .B2 (n_4511));
XOR2_X1 i_4604 (.Z (n_4497), .A (n_154), .B (n_4508));
XOR2_X1 i_4603 (.Z (n_4496), .A (n_4507), .B (n_4497));
NAND2_X1 i_4602 (.ZN (n_4495), .A1 (inputB[26]), .A2 (inputA[28]));
XOR2_X1 i_4601 (.Z (n_4494), .A (n_165), .B (n_4495));
AND2_X1 i_4600 (.ZN (n_4493), .A1 (inputB[28]), .A2 (inputA[26]));
NAND2_X1 i_4599 (.ZN (n_4492), .A1 (n_4494), .A2 (n_4493));
OAI21_X1 i_4598 (.ZN (n_4491), .A (n_4492), .B1 (n_4494), .B2 (n_4493));
OAI22_X1 i_4597 (.ZN (n_4490), .A1 (n_138), .A2 (n_137), .B1 (n_145), .B2 (n_139));
OAI21_X1 i_4596 (.ZN (n_4489), .A (n_4492), .B1 (n_165), .B2 (n_4495));
XOR2_X1 i_4595 (.Z (n_4488), .A (n_4490), .B (n_4489));
OAI21_X1 i_4594 (.ZN (n_4487), .A (n_147), .B1 (n_146), .B2 (n_140));
AOI22_X1 i_4593 (.ZN (n_4486), .A1 (n_4507), .A2 (n_4497), .B1 (n_4496), .B2 (n_4491));
XOR2_X1 i_4591 (.Z (n_4485), .A (n_4488), .B (n_4487));
NOR2_X1 i_4590 (.ZN (n_4484), .A1 (n_4486), .A2 (n_4485));
AOI21_X1 i_4589 (.ZN (n_4483), .A (n_4484), .B1 (n_4486), .B2 (n_4485));
AOI21_X1 i_4588 (.ZN (n_4482), .A (n_132), .B1 (n_4517), .B2 (n_133));
AOI21_X1 i_4587 (.ZN (n_4481), .A (n_4484), .B1 (n_4483), .B2 (n_4482));
INV_X1 i_4586 (.ZN (n_4480), .A (n_267));
INV_X1 i_4585 (.ZN (n_4478), .A (n_256));
INV_X1 i_4584 (.ZN (n_4477), .A (n_246));
INV_X1 i_4583 (.ZN (n_4476), .A (n_308));
INV_X1 i_4582 (.ZN (n_4475), .A (n_4388));
INV_X1 i_4581 (.ZN (n_4474), .A (n_175));
AOI22_X1 i_4580 (.ZN (n_4473), .A1 (n_425), .A2 (n_424), .B1 (n_423), .B2 (n_422));
AOI22_X1 i_4579 (.ZN (n_4472), .A1 (n_420), .A2 (n_419), .B1 (n_4480), .B2 (n_418));
AOI21_X1 i_4578 (.ZN (n_4471), .A (n_4404), .B1 (n_4402), .B2 (n_4396));
XNOR2_X1 i_4577 (.ZN (n_4470), .A (n_4472), .B (n_4471));
OAI22_X1 i_4576 (.ZN (n_4460), .A1 (n_4472), .A2 (n_4471), .B1 (n_4473), .B2 (n_4470));
XOR2_X1 i_4575 (.Z (n_4459), .A (n_228), .B (n_223));
NOR2_X1 i_4574 (.ZN (n_4458), .A1 (n_4460), .A2 (n_4459));
AOI21_X1 i_4573 (.ZN (n_4457), .A (n_4458), .B1 (n_4460), .B2 (n_4459));
NOR2_X1 i_4572 (.ZN (n_4456), .A1 (n_258), .A2 (n_4478));
XOR2_X1 i_4571 (.Z (n_4455), .A (n_255), .B (n_4456));
NOR2_X1 i_4570 (.ZN (n_4454), .A1 (n_254), .A2 (n_4477));
XOR2_X1 i_4569 (.Z (n_4453), .A (n_239), .B (n_4454));
NAND2_X1 i_4568 (.ZN (n_4452), .A1 (n_4455), .A2 (n_4453));
AOI22_X1 i_4567 (.ZN (n_4451), .A1 (n_4476), .A2 (n_307), .B1 (n_304), .B2 (n_303));
INV_X1 i_4566 (.ZN (n_4450), .A (n_4451));
NOR2_X1 i_4565 (.ZN (n_4449), .A1 (n_4455), .A2 (n_4453));
OAI21_X1 i_4564 (.ZN (n_4448), .A (n_4452), .B1 (n_4450), .B2 (n_4449));
AOI21_X1 i_4563 (.ZN (n_4447), .A (n_4458), .B1 (n_4457), .B2 (n_4448));
XOR2_X1 i_4562 (.Z (n_4446), .A (n_186), .B (n_185));
XOR2_X1 i_4561 (.Z (n_4445), .A (n_172), .B (n_171));
XOR2_X1 i_4559 (.Z (n_4444), .A (n_4446), .B (n_4445));
XNOR2_X1 i_4558 (.ZN (n_4443), .A (n_180), .B (n_179));
NAND2_X1 i_4557 (.ZN (n_4439), .A1 (n_4444), .A2 (n_4443));
OAI21_X1 i_4556 (.ZN (n_4438), .A (n_4439), .B1 (n_4446), .B2 (n_4445));
AOI22_X1 i_4555 (.ZN (n_4437), .A1 (n_4391), .A2 (n_4390), .B1 (n_4475), .B2 (n_4389));
NAND2_X1 i_4554 (.ZN (n_4436), .A1 (inputA[19]), .A2 (inputB[31]));
XOR2_X1 i_4553 (.Z (n_4435), .A (n_4474), .B (n_4436));
NOR2_X1 i_4552 (.ZN (n_4434), .A1 (n_481), .A2 (n_882));
AOI22_X1 i_4551 (.ZN (n_4433), .A1 (n_4474), .A2 (n_4436), .B1 (n_4435), .B2 (n_4434));
XNOR2_X1 i_4550 (.ZN (n_4432), .A (n_210), .B (n_209));
XOR2_X1 i_4549 (.Z (n_4431), .A (n_4433), .B (n_4432));
AOI22_X1 i_4548 (.ZN (n_4430), .A1 (n_4433), .A2 (n_4432), .B1 (n_4437), .B2 (n_4431));
XOR2_X1 i_4547 (.Z (n_4420), .A (n_4438), .B (n_4430));
XOR2_X1 i_4546 (.Z (n_4419), .A (n_4447), .B (n_4420));
NAND3_X1 i_4545 (.ZN (n_4418), .A1 (n_363), .A2 (inputA[29]), .A3 (inputB[21]));
OAI22_X1 i_4544 (.ZN (n_4417), .A1 (n_414), .A2 (n_123), .B1 (n_216), .B2 (n_122));
NAND2_X1 i_4543 (.ZN (n_4416), .A1 (n_4418), .A2 (n_4417));
XOR2_X1 i_4542 (.Z (n_4412), .A (n_373), .B (n_4416));
NOR2_X1 i_4541 (.ZN (n_4411), .A1 (n_275), .A2 (n_255));
AOI22_X1 i_4540 (.ZN (n_4410), .A1 (inputB[24]), .A2 (inputA[25]), .B1 (inputB[25]), .B2 (inputA[24]));
NOR2_X1 i_4539 (.ZN (n_4409), .A1 (n_4411), .A2 (n_4410));
XOR2_X1 i_4538 (.Z (n_4408), .A (n_257), .B (n_4409));
NOR2_X1 i_4537 (.ZN (n_4406), .A1 (n_4412), .A2 (n_4408));
AOI21_X1 i_4536 (.ZN (n_4405), .A (n_4406), .B1 (n_4412), .B2 (n_4408));
NOR2_X1 i_4535 (.ZN (n_4404), .A1 (n_329), .A2 (n_227));
AOI22_X1 i_4534 (.ZN (n_4403), .A1 (inputB[26]), .A2 (inputA[23]), .B1 (inputB[27]), .B2 (inputA[22]));
NOR2_X1 i_4533 (.ZN (n_4402), .A1 (n_4404), .A2 (n_4403));
NOR2_X1 i_4532 (.ZN (n_4396), .A1 (n_482), .A2 (n_127));
XNOR2_X1 i_4531 (.ZN (n_4392), .A (n_4402), .B (n_4396));
OAI21_X1 i_4530 (.ZN (n_4391), .A (n_4418), .B1 (n_373), .B2 (n_4416));
NAND2_X1 i_4529 (.ZN (n_4390), .A1 (inputB[19]), .A2 (inputA[31]));
XOR2_X1 i_4528 (.Z (n_4389), .A (n_4391), .B (n_4390));
AOI21_X1 i_4527 (.ZN (n_4388), .A (n_4411), .B1 (n_257), .B2 (n_4409));
AOI21_X1 i_4526 (.ZN (n_4387), .A (n_4406), .B1 (n_4405), .B2 (n_4392));
XNOR2_X1 i_4525 (.ZN (n_4386), .A (n_4389), .B (n_4388));
NOR2_X1 i_4524 (.ZN (n_4385), .A1 (n_4387), .A2 (n_4386));
AOI21_X1 i_4522 (.ZN (n_4384), .A (n_4385), .B1 (n_4387), .B2 (n_4386));
AOI22_X1 i_4521 (.ZN (n_4382), .A1 (n_261), .A2 (n_302), .B1 (n_269), .B2 (n_262));
INV_X1 i_4520 (.ZN (n_4381), .A (n_4382));
AOI21_X1 i_4519 (.ZN (n_4380), .A (n_4385), .B1 (n_4384), .B2 (n_4381));
INV_X1 i_4518 (.ZN (n_4379), .A (n_4028));
INV_X1 i_4517 (.ZN (n_4369), .A (n_3969));
INV_X1 i_4516 (.ZN (n_4368), .A (n_4010));
XNOR2_X1 i_4515 (.ZN (n_4367), .A (n_4132), .B (n_3984));
NAND2_X1 i_4514 (.ZN (n_4366), .A1 (inputB[7]), .A2 (inputA[31]));
OAI33_X1 i_4513 (.ZN (n_4365), .A1 (n_1131), .A2 (n_215), .A3 (n_4367), .B1 (n_3984)
    , .B2 (n_1127), .B3 (n_122));
XOR2_X1 i_4512 (.Z (n_4364), .A (n_4366), .B (n_4365));
NAND2_X1 i_4511 (.ZN (n_4354), .A1 (inputB[11]), .A2 (inputA[26]));
XNOR2_X1 i_4510 (.ZN (n_4353), .A (n_4134), .B (n_4354));
NAND2_X1 i_4509 (.ZN (n_4351), .A1 (inputB[13]), .A2 (inputA[24]));
OAI22_X1 i_4508 (.ZN (n_4350), .A1 (n_4134), .A2 (n_4354), .B1 (n_4353), .B2 (n_4351));
NAND2_X1 i_4507 (.ZN (n_4349), .A1 (inputB[17]), .A2 (inputA[19]));
NOR2_X1 i_4506 (.ZN (n_4347), .A1 (n_4033), .A2 (n_4349));
AOI22_X1 i_4505 (.ZN (n_4346), .A1 (inputB[18]), .A2 (inputA[19]), .B1 (inputB[17]), .B2 (inputA[20]));
NOR2_X1 i_4504 (.ZN (n_4345), .A1 (n_4347), .A2 (n_4346));
NAND2_X1 i_4503 (.ZN (n_4344), .A1 (inputB[19]), .A2 (inputA[18]));
INV_X1 i_4502 (.ZN (n_4342), .A (n_4344));
NOR2_X1 i_4501 (.ZN (n_4338), .A1 (n_4121), .A2 (n_3973));
AOI22_X1 i_4500 (.ZN (n_4337), .A1 (inputB[15]), .A2 (inputA[22]), .B1 (inputB[14]), .B2 (inputA[23]));
NOR2_X1 i_4499 (.ZN (n_4335), .A1 (n_4338), .A2 (n_4337));
NOR2_X1 i_4498 (.ZN (n_4334), .A1 (n_588), .A2 (n_482));
AOI21_X1 i_4497 (.ZN (n_4333), .A (n_4347), .B1 (n_4345), .B2 (n_4342));
AOI21_X1 i_4496 (.ZN (n_4332), .A (n_4338), .B1 (n_4335), .B2 (n_4334));
XNOR2_X1 i_4495 (.ZN (n_4321), .A (n_4333), .B (n_4332));
AOI22_X1 i_4494 (.ZN (n_4320), .A1 (inputB[22]), .A2 (inputA[15]), .B1 (inputB[21]), .B2 (inputA[16]));
AOI21_X1 i_4493 (.ZN (n_4319), .A (n_4320), .B1 (n_4153), .B2 (n_4027));
AOI22_X1 i_4492 (.ZN (n_4316), .A1 (n_4153), .A2 (n_4027), .B1 (n_4379), .B2 (n_4319));
OAI22_X1 i_4491 (.ZN (n_4315), .A1 (n_4333), .A2 (n_4332), .B1 (n_4321), .B2 (n_4316));
INV_X1 i_4490 (.ZN (n_4314), .A (n_4315));
AOI22_X1 i_4489 (.ZN (n_4313), .A1 (n_4366), .A2 (n_4365), .B1 (n_4364), .B2 (n_4350));
XOR2_X1 i_4488 (.Z (n_4312), .A (n_4314), .B (n_4313));
XOR2_X1 i_4487 (.Z (n_4311), .A (n_4200), .B (n_3983));
OAI21_X1 i_4486 (.ZN (n_4310), .A (n_4188), .B1 (n_4189), .B2 (n_4274));
INV_X1 i_4485 (.ZN (n_4309), .A (n_4310));
XOR2_X1 i_4484 (.Z (n_4308), .A (n_4179), .B (n_4237));
XOR2_X1 i_4483 (.Z (n_4303), .A (n_4309), .B (n_4308));
XNOR2_X1 i_4482 (.ZN (n_4302), .A (n_4171), .B (n_4170));
NAND2_X1 i_4480 (.ZN (n_4301), .A1 (n_4303), .A2 (n_4302));
OAI21_X1 i_4479 (.ZN (n_4300), .A (n_4301), .B1 (n_4309), .B2 (n_4308));
INV_X1 i_4478 (.ZN (n_4299), .A (n_4300));
AOI22_X1 i_4477 (.ZN (n_4298), .A1 (n_4314), .A2 (n_4313), .B1 (n_4312), .B2 (n_4311));
NOR2_X1 i_4476 (.ZN (n_4297), .A1 (n_4299), .A2 (n_4298));
AOI21_X1 i_4475 (.ZN (n_4296), .A (n_4297), .B1 (n_4299), .B2 (n_4298));
OAI22_X1 i_4474 (.ZN (n_4295), .A1 (n_3985), .A2 (n_3978), .B1 (n_4369), .B2 (n_3977));
AOI21_X1 i_4473 (.ZN (n_4294), .A (n_4095), .B1 (n_4093), .B2 (n_4091));
XNOR2_X1 i_4472 (.ZN (n_4293), .A (n_4295), .B (n_4294));
AOI22_X1 i_4471 (.ZN (n_4292), .A1 (n_4368), .A2 (n_4029), .B1 (n_4009), .B2 (n_3993));
XOR2_X1 i_4470 (.Z (n_4291), .A (n_4293), .B (n_4292));
AOI21_X1 i_4469 (.ZN (n_4290), .A (n_4297), .B1 (n_4296), .B2 (n_4291));
XNOR2_X1 i_4468 (.ZN (n_4289), .A (n_3860), .B (n_3859));
OAI21_X1 i_4467 (.ZN (n_4288), .A (n_3802), .B1 (n_3803), .B2 (n_3622));
XOR2_X1 i_4466 (.Z (n_4287), .A (n_4289), .B (n_4288));
XOR2_X1 i_4465 (.Z (n_4286), .A (n_3785), .B (n_3784));
XOR2_X1 i_4464 (.Z (n_4285), .A (n_3745), .B (n_3739));
NAND2_X1 i_4463 (.ZN (n_4284), .A1 (n_3733), .A2 (n_3735));
XNOR2_X1 i_4462 (.ZN (n_4282), .A (n_3731), .B (n_4284));
NOR2_X1 i_4461 (.ZN (n_4281), .A1 (n_4226), .A2 (n_4225));
XOR2_X1 i_4460 (.Z (n_4280), .A (n_4222), .B (n_4281));
XOR2_X1 i_4459 (.Z (n_4279), .A (n_4282), .B (n_4280));
XNOR2_X1 i_4458 (.ZN (n_4278), .A (n_4287), .B (n_4286));
XOR2_X1 i_4457 (.Z (n_4277), .A (n_4285), .B (n_4279));
XOR2_X1 i_4456 (.Z (n_4276), .A (n_4278), .B (n_4277));
AOI22_X1 i_4455 (.ZN (n_4275), .A1 (n_4278), .A2 (n_4277), .B1 (n_4290), .B2 (n_4276));
INV_X1 i_4454 (.ZN (n_4274), .A (n_3992));
OR2_X1 i_4453 (.ZN (n_4273), .A1 (n_3718), .A2 (n_3784));
AOI22_X1 i_4452 (.ZN (n_4272), .A1 (inputA[18]), .A2 (inputB[22]), .B1 (inputA[19]), .B2 (inputB[21]));
INV_X1 i_4451 (.ZN (n_4271), .A (n_4272));
NAND2_X1 i_4450 (.ZN (n_4261), .A1 (n_4273), .A2 (n_4271));
AND2_X1 i_4449 (.ZN (n_4260), .A1 (inputA[23]), .A2 (inputB[17]));
XOR2_X1 i_4448 (.Z (n_4259), .A (n_3820), .B (n_4260));
OAI21_X1 i_4447 (.ZN (n_4258), .A (n_4273), .B1 (n_3788), .B2 (n_4261));
OAI33_X1 i_4446 (.ZN (n_4257), .A1 (n_314), .A2 (n_482), .A3 (n_4259), .B1 (n_3820)
    , .B2 (n_881), .B3 (n_213));
XOR2_X1 i_4445 (.Z (n_4256), .A (n_4258), .B (n_4257));
NOR2_X1 i_4444 (.ZN (n_4255), .A1 (n_3680), .A2 (n_3597));
AOI22_X1 i_4443 (.ZN (n_4254), .A1 (inputA[17]), .A2 (inputB[23]), .B1 (inputA[16]), .B2 (inputB[24]));
NOR2_X1 i_4442 (.ZN (n_4248), .A1 (n_4255), .A2 (n_4254));
OAI22_X1 i_4441 (.ZN (n_4246), .A1 (n_3680), .A2 (n_3597), .B1 (n_3689), .B2 (n_4254));
INV_X1 i_4440 (.ZN (n_4245), .A (n_4246));
AOI22_X1 i_4439 (.ZN (n_4244), .A1 (n_4258), .A2 (n_4257), .B1 (n_4256), .B2 (n_4246));
NAND2_X1 i_4438 (.ZN (n_4243), .A1 (inputA[28]), .A2 (inputB[12]));
XNOR2_X1 i_4437 (.ZN (n_4242), .A (n_3858), .B (n_4243));
NAND2_X1 i_4436 (.ZN (n_4241), .A1 (inputA[27]), .A2 (inputB[13]));
NAND2_X1 i_4435 (.ZN (n_4240), .A1 (inputA[31]), .A2 (inputB[10]));
OAI22_X1 i_4434 (.ZN (n_4239), .A1 (n_3858), .A2 (n_4243), .B1 (n_4242), .B2 (n_4241));
XOR2_X1 i_4433 (.Z (n_4238), .A (n_4240), .B (n_4239));
NOR2_X1 i_4432 (.ZN (n_4237), .A1 (n_586), .A2 (n_483));
NAND3_X1 i_4431 (.ZN (n_4236), .A1 (inputB[15]), .A2 (n_4237), .A3 (inputA[26]));
OAI22_X1 i_4430 (.ZN (n_4235), .A1 (n_586), .A2 (n_214), .B1 (n_483), .B2 (n_587));
NAND2_X1 i_4429 (.ZN (n_4234), .A1 (n_4236), .A2 (n_4235));
NAND2_X1 i_4428 (.ZN (n_4233), .A1 (inputA[24]), .A2 (inputB[16]));
OAI21_X1 i_4426 (.ZN (n_4232), .A (n_4236), .B1 (n_4234), .B2 (n_4233));
AOI22_X1 i_4425 (.ZN (n_4227), .A1 (n_4240), .A2 (n_4239), .B1 (n_4238), .B2 (n_4232));
NOR2_X1 i_4424 (.ZN (n_4226), .A1 (n_3638), .A2 (n_3584));
AOI22_X1 i_4423 (.ZN (n_4225), .A1 (inputA[11]), .A2 (inputB[30]), .B1 (inputA[12]), .B2 (inputB[29]));
INV_X1 i_4422 (.ZN (n_4224), .A (n_4225));
NAND2_X1 i_4421 (.ZN (n_4222), .A1 (inputA[10]), .A2 (inputB[31]));
AOI21_X1 i_4420 (.ZN (n_4221), .A (n_4226), .B1 (n_4224), .B2 (n_4222));
XNOR2_X1 i_4419 (.ZN (n_4220), .A (n_4227), .B (n_4221));
XNOR2_X1 i_4418 (.ZN (n_4218), .A (n_4244), .B (n_4220));
NOR2_X1 i_4417 (.ZN (n_4217), .A1 (n_1131), .A2 (n_123));
NAND2_X1 i_4416 (.ZN (n_4216), .A1 (inputA[31]), .A2 (inputB[8]));
NAND2_X1 i_4415 (.ZN (n_4215), .A1 (n_4217), .A2 (n_4216));
NOR2_X1 i_4414 (.ZN (n_4214), .A1 (n_4217), .A2 (n_4216));
AOI21_X1 i_4413 (.ZN (n_4200), .A (n_4214), .B1 (n_4217), .B2 (n_4216));
NAND2_X1 i_4412 (.ZN (n_4199), .A1 (inputA[31]), .A2 (inputB[9]));
OAI21_X1 i_4411 (.ZN (n_4198), .A (n_4215), .B1 (n_3983), .B2 (n_4214));
XOR2_X1 i_4410 (.Z (n_4197), .A (n_4199), .B (n_4198));
NOR2_X1 i_4409 (.ZN (n_4196), .A1 (n_1131), .A2 (n_124));
AOI22_X1 i_4408 (.ZN (n_4195), .A1 (n_4199), .A2 (n_4198), .B1 (n_4197), .B2 (n_4196));
XNOR2_X1 i_4407 (.ZN (n_4194), .A (n_3854), .B (n_3853));
NAND2_X1 i_4406 (.ZN (n_4193), .A1 (n_4195), .A2 (n_4194));
OAI21_X1 i_4405 (.ZN (n_4192), .A (n_4193), .B1 (n_4195), .B2 (n_4194));
NOR2_X1 i_4404 (.ZN (n_4191), .A1 (n_3987), .A2 (n_4243));
AOI22_X1 i_4403 (.ZN (n_4190), .A1 (inputA[28]), .A2 (inputB[11]), .B1 (inputA[27]), .B2 (inputB[12]));
NOR2_X1 i_4402 (.ZN (n_4189), .A1 (n_4191), .A2 (n_4190));
NAND2_X1 i_4401 (.ZN (n_4188), .A1 (n_4274), .A2 (n_4189));
NOR2_X1 i_4400 (.ZN (n_4187), .A1 (n_3973), .A2 (n_4233));
AOI22_X1 i_4399 (.ZN (n_4180), .A1 (inputA[23]), .A2 (inputB[16]), .B1 (inputA[24]), .B2 (inputB[15]));
NOR2_X1 i_4398 (.ZN (n_4179), .A1 (n_4187), .A2 (n_4180));
AOI21_X1 i_4397 (.ZN (n_4178), .A (n_4191), .B1 (n_4274), .B2 (n_4189));
AOI21_X1 i_4396 (.ZN (n_4177), .A (n_4187), .B1 (n_4237), .B2 (n_4179));
NOR2_X1 i_4395 (.ZN (n_4176), .A1 (n_4178), .A2 (n_4177));
AOI21_X1 i_4394 (.ZN (n_4175), .A (n_4176), .B1 (n_4178), .B2 (n_4177));
OR2_X1 i_4393 (.ZN (n_4174), .A1 (n_3820), .A2 (n_4032));
AOI22_X1 i_4392 (.ZN (n_4173), .A1 (inputA[22]), .A2 (inputB[17]), .B1 (inputA[21]), .B2 (inputB[18]));
INV_X1 i_4391 (.ZN (n_4172), .A (n_4173));
NAND2_X1 i_4390 (.ZN (n_4171), .A1 (n_4174), .A2 (n_4172));
NAND2_X1 i_4389 (.ZN (n_4170), .A1 (inputA[20]), .A2 (inputB[19]));
OAI21_X1 i_4388 (.ZN (n_4169), .A (n_4174), .B1 (n_4171), .B2 (n_4170));
AOI21_X1 i_4387 (.ZN (n_4168), .A (n_4176), .B1 (n_4175), .B2 (n_4169));
INV_X1 i_4386 (.ZN (n_4167), .A (n_4168));
OAI21_X1 i_4385 (.ZN (n_4165), .A (n_4193), .B1 (n_4192), .B2 (n_4167));
XOR2_X1 i_4384 (.Z (n_4164), .A (n_4218), .B (n_4165));
INV_X1 i_4383 (.ZN (n_4163), .A (n_4349));
INV_X1 i_4382 (.ZN (n_4162), .A (inputA[10]));
NOR2_X1 i_4380 (.ZN (n_4161), .A1 (n_654), .A2 (n_4344));
NOR2_X1 i_4379 (.ZN (n_4160), .A1 (n_50), .A2 (n_4161));
NAND2_X1 i_4378 (.ZN (n_4159), .A1 (n_4163), .A2 (n_4160));
NAND2_X1 i_4377 (.ZN (n_4158), .A1 (inputA[13]), .A2 (inputB[23]));
XNOR2_X1 i_4376 (.ZN (n_4157), .A (n_1047), .B (n_4158));
OAI21_X1 i_4375 (.ZN (n_4156), .A (n_4159), .B1 (n_654), .B2 (n_4344));
OAI33_X1 i_4374 (.ZN (n_4155), .A1 (n_1136), .A2 (n_219), .A3 (n_4157), .B1 (n_667)
    , .B2 (n_461), .B3 (n_4158));
XOR2_X1 i_4373 (.Z (n_4154), .A (n_4156), .B (n_4155));
NOR2_X1 i_4372 (.ZN (n_4153), .A1 (n_478), .A2 (n_216));
NOR2_X1 i_4371 (.ZN (n_4152), .A1 (n_865), .A2 (n_414));
NAND2_X1 i_4370 (.ZN (n_4151), .A1 (n_4153), .A2 (n_4152));
OAI21_X1 i_4369 (.ZN (n_4150), .A (n_4151), .B1 (n_4153), .B2 (n_4152));
NAND2_X1 i_4368 (.ZN (n_4149), .A1 (inputA[14]), .A2 (inputB[22]));
OAI21_X1 i_4367 (.ZN (n_4136), .A (n_4151), .B1 (n_4150), .B2 (n_4149));
NAND2_X1 i_4366 (.ZN (n_4135), .A1 (n_48), .A2 (n_49));
NAND2_X1 i_4365 (.ZN (n_4134), .A1 (inputA[25]), .A2 (inputB[12]));
NOR2_X1 i_4364 (.ZN (n_4133), .A1 (n_1015), .A2 (n_4134));
NAND2_X1 i_4363 (.ZN (n_4132), .A1 (inputA[28]), .A2 (inputB[9]));
NOR3_X1 i_4362 (.ZN (n_4131), .A1 (n_669), .A2 (n_4132), .A3 (n_215));
AOI22_X1 i_4361 (.ZN (n_4130), .A1 (inputA[28]), .A2 (inputB[8]), .B1 (inputA[27]), .B2 (inputB[9]));
NOR2_X1 i_4360 (.ZN (n_4129), .A1 (n_4131), .A2 (n_4130));
NOR2_X1 i_4359 (.ZN (n_4128), .A1 (n_1131), .A2 (n_214));
OAI21_X1 i_4358 (.ZN (n_4127), .A (n_4135), .B1 (n_1015), .B2 (n_4134));
AOI21_X1 i_4357 (.ZN (n_4126), .A (n_4131), .B1 (n_4129), .B2 (n_4128));
INV_X1 i_4356 (.ZN (n_4125), .A (n_4126));
NAND2_X1 i_4355 (.ZN (n_4124), .A1 (n_4127), .A2 (n_4125));
OAI21_X1 i_4354 (.ZN (n_4123), .A (n_4124), .B1 (n_4127), .B2 (n_4125));
NAND2_X1 i_4353 (.ZN (n_4121), .A1 (inputA[22]), .A2 (inputB[14]));
NOR2_X1 i_4352 (.ZN (n_4120), .A1 (n_1028), .A2 (n_4121));
AOI21_X1 i_4351 (.ZN (n_4119), .A (n_4120), .B1 (n_1028), .B2 (n_4121));
NOR2_X1 i_4350 (.ZN (n_4118), .A1 (n_588), .A2 (n_481));
AOI21_X1 i_4349 (.ZN (n_4117), .A (n_4120), .B1 (n_4119), .B2 (n_4118));
AOI22_X1 i_4348 (.ZN (n_4116), .A1 (n_4156), .A2 (n_4155), .B1 (n_4154), .B2 (n_4136));
OAI21_X1 i_4347 (.ZN (n_4115), .A (n_4124), .B1 (n_4123), .B2 (n_4117));
INV_X1 i_4346 (.ZN (n_4114), .A (n_4115));
NOR2_X1 i_4345 (.ZN (n_4113), .A1 (n_4116), .A2 (n_4114));
AOI21_X1 i_4344 (.ZN (n_4112), .A (n_4113), .B1 (n_4116), .B2 (n_4114));
NOR2_X1 i_4343 (.ZN (n_4111), .A1 (n_879), .A2 (n_123));
NAND2_X1 i_4342 (.ZN (n_4110), .A1 (inputA[31]), .A2 (inputB[5]));
XOR2_X1 i_4341 (.Z (n_4109), .A (n_4111), .B (n_4110));
NOR2_X1 i_4340 (.ZN (n_4108), .A1 (n_878), .A2 (n_125));
AOI22_X1 i_4339 (.ZN (n_4107), .A1 (n_4111), .A2 (n_4110), .B1 (n_756), .B2 (n_4109));
XNOR2_X1 i_4338 (.ZN (n_4099), .A (n_4108), .B (n_4107));
NAND2_X1 i_4337 (.ZN (n_4098), .A1 (inputA[30]), .A2 (inputB[7]));
OAI22_X1 i_4336 (.ZN (n_4097), .A1 (n_4108), .A2 (n_4107), .B1 (n_4099), .B2 (n_4098));
NAND2_X1 i_4335 (.ZN (n_4096), .A1 (inputA[9]), .A2 (inputB[29]));
NOR2_X1 i_4334 (.ZN (n_4095), .A1 (n_3631), .A2 (n_4096));
AOI22_X1 i_4333 (.ZN (n_4094), .A1 (inputA[9]), .A2 (inputB[30]), .B1 (inputA[10]), .B2 (inputB[29]));
NOR2_X1 i_4332 (.ZN (n_4093), .A1 (n_4095), .A2 (n_4094));
NAND2_X1 i_4331 (.ZN (n_4091), .A1 (inputA[8]), .A2 (inputB[31]));
AOI21_X1 i_4330 (.ZN (n_4090), .A (n_4113), .B1 (n_4112), .B2 (n_4097));
INV_X1 i_4329 (.ZN (n_4089), .A (n_4090));
XOR2_X1 i_4328 (.Z (n_4088), .A (n_4093), .B (n_4091));
XOR2_X1 i_4327 (.Z (n_4086), .A (n_4089), .B (n_4088));
NOR2_X1 i_4326 (.ZN (n_4083), .A1 (n_864), .A2 (n_129));
XNOR2_X1 i_4325 (.ZN (n_4082), .A (n_4096), .B (n_4083));
NAND2_X1 i_4324 (.ZN (n_4067), .A1 (inputA[8]), .A2 (inputB[30]));
AND2_X1 i_4323 (.ZN (n_4066), .A1 (inputA[11]), .A2 (inputB[27]));
XOR2_X1 i_4322 (.Z (n_4065), .A (n_3676), .B (n_4066));
NOR2_X1 i_4321 (.ZN (n_4064), .A1 (n_129), .A2 (n_1349));
NAND2_X1 i_4320 (.ZN (n_4063), .A1 (inputA[8]), .A2 (inputB[29]));
XNOR2_X1 i_4319 (.ZN (n_4062), .A (n_4064), .B (n_4063));
OAI33_X1 i_4317 (.ZN (n_4061), .A1 (n_864), .A2 (n_882), .A3 (n_4062), .B1 (n_1551)
    , .B2 (n_128), .B3 (n_4064));
NAND2_X1 i_4316 (.ZN (n_4060), .A1 (inputA[10]), .A2 (inputB[27]));
NAND2_X1 i_4315 (.ZN (n_4059), .A1 (inputA[11]), .A2 (inputB[26]));
XNOR2_X1 i_4314 (.ZN (n_4058), .A (n_4060), .B (n_4059));
NAND2_X1 i_4313 (.ZN (n_4057), .A1 (inputA[9]), .A2 (inputB[28]));
NOR2_X1 i_4312 (.ZN (n_4053), .A1 (n_3697), .A2 (n_4158));
AOI22_X1 i_4311 (.ZN (n_4052), .A1 (inputA[14]), .A2 (inputB[23]), .B1 (inputA[13]), .B2 (inputB[24]));
NOR2_X1 i_4310 (.ZN (n_4051), .A1 (n_4053), .A2 (n_4052));
NOR2_X1 i_4309 (.ZN (n_4050), .A1 (n_219), .A2 (n_667));
AOI21_X1 i_4308 (.ZN (n_4049), .A (n_4053), .B1 (n_4051), .B2 (n_4050));
OAI22_X1 i_4307 (.ZN (n_4046), .A1 (n_4060), .A2 (n_4059), .B1 (n_4058), .B2 (n_4057));
INV_X1 i_4306 (.ZN (n_4045), .A (n_4046));
NOR2_X1 i_4305 (.ZN (n_4044), .A1 (n_4049), .A2 (n_4045));
AOI21_X1 i_4304 (.ZN (n_4042), .A (n_4044), .B1 (n_4049), .B2 (n_4045));
OAI33_X1 i_4303 (.ZN (n_4041), .A1 (n_4162), .A2 (n_127), .A3 (n_4065), .B1 (n_667)
    , .B2 (n_126), .B3 (n_4059));
OAI22_X1 i_4302 (.ZN (n_4040), .A1 (n_4096), .A2 (n_4083), .B1 (n_4082), .B2 (n_4067));
XNOR2_X1 i_4301 (.ZN (n_4039), .A (n_4041), .B (n_4040));
AOI21_X1 i_4300 (.ZN (n_4037), .A (n_4044), .B1 (n_4061), .B2 (n_4042));
NOR2_X1 i_4299 (.ZN (n_4036), .A1 (n_4039), .A2 (n_4037));
AOI21_X1 i_4298 (.ZN (n_4035), .A (n_4036), .B1 (n_4039), .B2 (n_4037));
AOI22_X1 i_4297 (.ZN (n_4034), .A1 (n_4089), .A2 (n_4088), .B1 (n_4086), .B2 (n_4035));
NAND2_X1 i_4296 (.ZN (n_4033), .A1 (inputA[20]), .A2 (inputB[18]));
NAND2_X1 i_4295 (.ZN (n_4032), .A1 (inputA[21]), .A2 (inputB[17]));
XNOR2_X1 i_4294 (.ZN (n_4031), .A (n_4033), .B (n_4032));
NAND2_X1 i_4293 (.ZN (n_4030), .A1 (inputA[19]), .A2 (inputB[19]));
OAI22_X1 i_4292 (.ZN (n_4029), .A1 (n_4033), .A2 (n_4032), .B1 (n_4031), .B2 (n_4030));
NAND2_X1 i_4291 (.ZN (n_4028), .A1 (inputA[17]), .A2 (inputB[20]));
NOR2_X1 i_4290 (.ZN (n_4027), .A1 (n_865), .A2 (n_217));
NOR2_X1 i_4289 (.ZN (n_4026), .A1 (n_3718), .A2 (n_4028));
AOI22_X1 i_4288 (.ZN (n_4025), .A1 (inputA[18]), .A2 (inputB[20]), .B1 (inputA[17]), .B2 (inputB[21]));
NOR2_X1 i_4287 (.ZN (n_4024), .A1 (n_4026), .A2 (n_4025));
AOI21_X1 i_4286 (.ZN (n_4010), .A (n_4026), .B1 (n_4027), .B2 (n_4024));
XNOR2_X1 i_4285 (.ZN (n_4009), .A (n_4029), .B (n_4010));
NAND2_X1 i_4284 (.ZN (n_4008), .A1 (inputA[15]), .A2 (inputB[23]));
XNOR2_X1 i_4283 (.ZN (n_4007), .A (n_3697), .B (n_4008));
NAND2_X1 i_4282 (.ZN (n_4006), .A1 (inputA[13]), .A2 (inputB[25]));
OAI22_X1 i_4281 (.ZN (n_3993), .A1 (n_3697), .A2 (n_4008), .B1 (n_4007), .B2 (n_4006));
NAND2_X1 i_4280 (.ZN (n_3992), .A1 (inputA[26]), .A2 (inputB[13]));
NOR2_X1 i_4279 (.ZN (n_3991), .A1 (n_4134), .A2 (n_3992));
INV_X1 i_4278 (.ZN (n_3990), .A (n_3991));
AOI22_X1 i_4277 (.ZN (n_3989), .A1 (inputA[25]), .A2 (inputB[13]), .B1 (inputA[26]), .B2 (inputB[12]));
NOR2_X1 i_4276 (.ZN (n_3988), .A1 (n_3991), .A2 (n_3989));
NAND2_X1 i_4275 (.ZN (n_3987), .A1 (inputA[27]), .A2 (inputB[11]));
AOI21_X1 i_4274 (.ZN (n_3986), .A (n_3989), .B1 (n_3990), .B2 (n_3987));
INV_X1 i_4273 (.ZN (n_3985), .A (n_3986));
NAND2_X1 i_4272 (.ZN (n_3984), .A1 (inputA[29]), .A2 (inputB[8]));
NAND2_X1 i_4271 (.ZN (n_3983), .A1 (inputA[30]), .A2 (inputB[9]));
NOR2_X1 i_4270 (.ZN (n_3982), .A1 (n_3984), .A2 (n_3983));
AOI22_X1 i_4269 (.ZN (n_3981), .A1 (inputA[30]), .A2 (inputB[8]), .B1 (inputA[29]), .B2 (inputB[9]));
NOR2_X1 i_4268 (.ZN (n_3980), .A1 (n_3982), .A2 (n_3981));
NOR2_X1 i_4267 (.ZN (n_3979), .A1 (n_1131), .A2 (n_122));
AOI21_X1 i_4266 (.ZN (n_3978), .A (n_3982), .B1 (n_3980), .B2 (n_3979));
XOR2_X1 i_4265 (.Z (n_3977), .A (n_3986), .B (n_3978));
NAND2_X1 i_4264 (.ZN (n_3973), .A1 (inputA[23]), .A2 (inputB[15]));
NAND2_X1 i_4263 (.ZN (n_3972), .A1 (inputA[24]), .A2 (inputB[14]));
XNOR2_X1 i_4262 (.ZN (n_3971), .A (n_3973), .B (n_3972));
NAND2_X1 i_4261 (.ZN (n_3970), .A1 (inputA[22]), .A2 (inputB[16]));
OAI22_X1 i_4260 (.ZN (n_3969), .A1 (n_3973), .A2 (n_3972), .B1 (n_3971), .B2 (n_3970));
XOR2_X1 i_4259 (.Z (n_3967), .A (n_4009), .B (n_3993));
XNOR2_X1 i_4258 (.ZN (n_3966), .A (n_3977), .B (n_3969));
XOR2_X1 i_4256 (.Z (n_3965), .A (n_3967), .B (n_3966));
XOR2_X1 i_4255 (.Z (n_3964), .A (n_4027), .B (n_4024));
XOR2_X1 i_4254 (.Z (n_3963), .A (n_4031), .B (n_4030));
NOR2_X1 i_4253 (.ZN (n_3962), .A1 (n_3964), .A2 (n_3963));
AOI21_X1 i_4252 (.ZN (n_3961), .A (n_3962), .B1 (n_3964), .B2 (n_3963));
XNOR2_X1 i_4251 (.ZN (n_3960), .A (n_4007), .B (n_4006));
AOI21_X1 i_4250 (.ZN (n_3959), .A (n_3962), .B1 (n_3961), .B2 (n_3960));
XOR2_X1 i_4249 (.Z (n_3951), .A (n_3640), .B (n_3639));
XNOR2_X1 i_4248 (.ZN (n_3950), .A (n_3631), .B (n_3636));
XOR2_X1 i_4247 (.Z (n_3949), .A (n_3951), .B (n_3950));
AOI21_X1 i_4246 (.ZN (n_3948), .A (n_4036), .B1 (n_4041), .B2 (n_4040));
AOI22_X1 i_4245 (.ZN (n_3947), .A1 (n_3967), .A2 (n_3966), .B1 (n_3965), .B2 (n_3959));
XOR2_X1 i_4244 (.Z (n_3946), .A (n_3949), .B (n_3948));
XOR2_X1 i_4243 (.Z (n_3945), .A (n_3947), .B (n_3946));
AOI22_X1 i_4242 (.ZN (n_3944), .A1 (n_3947), .A2 (n_3946), .B1 (n_4034), .B2 (n_3945));
OR2_X1 i_4241 (.ZN (n_3941), .A1 (n_671), .A2 (n_123));
NAND2_X1 i_4240 (.ZN (n_3940), .A1 (inputB[12]), .A2 (inputA[30]));
AND2_X1 i_4239 (.ZN (n_3939), .A1 (inputB[11]), .A2 (inputA[31]));
XNOR2_X1 i_4238 (.ZN (n_3938), .A (n_3940), .B (n_3939));
XOR2_X1 i_4237 (.Z (n_3937), .A (n_3941), .B (n_3938));
XNOR2_X1 i_4236 (.ZN (n_3909), .A (n_3618), .B (n_3613));
NOR2_X1 i_4235 (.ZN (n_3908), .A1 (n_3937), .A2 (n_3909));
AOI21_X1 i_4234 (.ZN (n_3907), .A (n_3908), .B1 (n_3937), .B2 (n_3909));
NAND2_X1 i_4233 (.ZN (n_3906), .A1 (inputB[16]), .A2 (inputA[26]));
XNOR2_X1 i_4232 (.ZN (n_3897), .A (n_3623), .B (n_3906));
AOI21_X1 i_4231 (.ZN (n_3896), .A (n_3908), .B1 (n_3907), .B2 (n_3897));
XOR2_X1 i_4230 (.Z (n_3895), .A (n_3593), .B (n_3592));
XOR2_X1 i_4229 (.Z (n_3894), .A (n_3607), .B (n_3606));
NOR2_X1 i_4228 (.ZN (n_3892), .A1 (n_3895), .A2 (n_3894));
AOI21_X1 i_4227 (.ZN (n_3891), .A (n_3892), .B1 (n_3895), .B2 (n_3894));
XNOR2_X1 i_4226 (.ZN (n_3890), .A (n_3601), .B (n_3598));
AOI21_X1 i_4225 (.ZN (n_3889), .A (n_3892), .B1 (n_3891), .B2 (n_3890));
XOR2_X1 i_4224 (.Z (n_3888), .A (n_3896), .B (n_3889));
OAI22_X1 i_4223 (.ZN (n_3871), .A1 (n_3736), .A2 (n_3725), .B1 (n_3782), .B2 (n_3737));
OR3_X1 i_4222 (.ZN (n_3862), .A1 (n_3625), .A2 (n_214), .A3 (n_586));
OAI22_X1 i_4221 (.ZN (n_3861), .A1 (n_586), .A2 (n_215), .B1 (n_214), .B2 (n_587));
NAND2_X1 i_4220 (.ZN (n_3860), .A1 (n_3862), .A2 (n_3861));
NAND2_X1 i_4219 (.ZN (n_3859), .A1 (inputB[16]), .A2 (inputA[25]));
NAND2_X1 i_4218 (.ZN (n_3858), .A1 (inputB[11]), .A2 (inputA[29]));
AOI22_X1 i_4217 (.ZN (n_3856), .A1 (inputB[11]), .A2 (inputA[30]), .B1 (inputB[12]), .B2 (inputA[29]));
INV_X1 i_4216 (.ZN (n_3855), .A (n_3856));
OAI21_X1 i_4215 (.ZN (n_3854), .A (n_3855), .B1 (n_3940), .B2 (n_3858));
NAND2_X1 i_4214 (.ZN (n_3853), .A1 (inputB[13]), .A2 (inputA[28]));
OAI21_X1 i_4213 (.ZN (n_3852), .A (n_3862), .B1 (n_3860), .B2 (n_3859));
OAI22_X1 i_4212 (.ZN (n_3823), .A1 (n_3940), .A2 (n_3858), .B1 (n_3854), .B2 (n_3853));
NAND2_X1 i_4211 (.ZN (n_3822), .A1 (n_3852), .A2 (n_3823));
OAI21_X1 i_4210 (.ZN (n_3821), .A (n_3822), .B1 (n_3852), .B2 (n_3823));
NAND2_X1 i_4209 (.ZN (n_3820), .A1 (inputB[18]), .A2 (inputA[22]));
NOR2_X1 i_4208 (.ZN (n_3817), .A1 (n_3613), .A2 (n_3820));
AOI22_X1 i_4207 (.ZN (n_3816), .A1 (inputB[18]), .A2 (inputA[23]), .B1 (inputB[19]), .B2 (inputA[22]));
NOR2_X1 i_4206 (.ZN (n_3803), .A1 (n_3817), .A2 (n_3816));
NAND2_X1 i_4205 (.ZN (n_3802), .A1 (n_3622), .A2 (n_3803));
AOI21_X1 i_4204 (.ZN (n_3801), .A (n_3817), .B1 (n_3622), .B2 (n_3803));
OAI21_X1 i_4203 (.ZN (n_3800), .A (n_3822), .B1 (n_3821), .B2 (n_3801));
XOR2_X1 i_4202 (.Z (n_3799), .A (n_3871), .B (n_3800));
OAI22_X1 i_4201 (.ZN (n_3797), .A1 (n_3940), .A2 (n_3939), .B1 (n_3941), .B2 (n_3938));
NAND2_X1 i_4199 (.ZN (n_3795), .A1 (inputB[12]), .A2 (inputA[31]));
XOR2_X1 i_4198 (.Z (n_3794), .A (n_3797), .B (n_3795));
NOR2_X1 i_4197 (.ZN (n_3793), .A1 (n_671), .A2 (n_124));
XOR2_X1 i_4196 (.Z (n_3791), .A (n_3794), .B (n_3793));
XOR2_X1 i_4195 (.Z (n_3790), .A (n_3799), .B (n_3791));
XOR2_X1 i_4194 (.Z (n_3789), .A (n_3888), .B (n_3790));
NAND2_X1 i_4193 (.ZN (n_3788), .A1 (inputA[20]), .A2 (inputB[20]));
NOR2_X1 i_4191 (.ZN (n_3787), .A1 (n_3609), .A2 (n_3788));
AOI22_X1 i_4190 (.ZN (n_3786), .A1 (inputA[20]), .A2 (inputB[21]), .B1 (inputA[21]), .B2 (inputB[20]));
NOR2_X1 i_4189 (.ZN (n_3785), .A1 (n_3787), .A2 (n_3786));
NAND2_X1 i_4188 (.ZN (n_3784), .A1 (inputA[19]), .A2 (inputB[22]));
INV_X1 i_4187 (.ZN (n_3783), .A (n_3784));
AOI21_X1 i_4186 (.ZN (n_3782), .A (n_3787), .B1 (n_3785), .B2 (n_3783));
NAND2_X1 i_4185 (.ZN (n_3777), .A1 (inputA[14]), .A2 (inputB[26]));
NOR2_X1 i_4184 (.ZN (n_3776), .A1 (n_3603), .A2 (n_3777));
AOI22_X1 i_4183 (.ZN (n_3775), .A1 (inputA[14]), .A2 (inputB[27]), .B1 (inputA[15]), .B2 (inputB[26]));
NOR2_X1 i_4182 (.ZN (n_3745), .A1 (n_3776), .A2 (n_3775));
NOR2_X1 i_4181 (.ZN (n_3739), .A1 (n_529), .A2 (n_127));
AOI21_X1 i_4180 (.ZN (n_3737), .A (n_3776), .B1 (n_3745), .B2 (n_3739));
XNOR2_X1 i_4179 (.ZN (n_3736), .A (n_3782), .B (n_3737));
OAI21_X1 i_4178 (.ZN (n_3735), .A (n_3597), .B1 (n_479), .B2 (n_218));
NOR3_X1 i_4177 (.ZN (n_3734), .A1 (n_3597), .A2 (n_479), .A3 (n_218));
INV_X1 i_4176 (.ZN (n_3733), .A (n_3734));
NOR2_X1 i_4175 (.ZN (n_3731), .A1 (n_865), .A2 (n_219));
OAI21_X1 i_4174 (.ZN (n_3725), .A (n_3735), .B1 (n_3734), .B2 (n_3731));
XOR2_X1 i_4173 (.Z (n_3724), .A (n_3585), .B (n_3584));
XOR2_X1 i_4172 (.Z (n_3723), .A (n_3736), .B (n_3725));
NOR2_X1 i_4171 (.ZN (n_3722), .A1 (n_3724), .A2 (n_3723));
AOI21_X1 i_4170 (.ZN (n_3721), .A (n_3722), .B1 (n_3724), .B2 (n_3723));
NAND2_X1 i_4169 (.ZN (n_3718), .A1 (inputA[18]), .A2 (inputB[21]));
NAND2_X1 i_4168 (.ZN (n_3717), .A1 (inputA[19]), .A2 (inputB[20]));
XNOR2_X1 i_4167 (.ZN (n_3716), .A (n_3718), .B (n_3717));
NAND2_X1 i_4166 (.ZN (n_3715), .A1 (inputA[17]), .A2 (inputB[22]));
NAND2_X1 i_4165 (.ZN (n_3697), .A1 (inputA[14]), .A2 (inputB[24]));
NAND2_X1 i_4164 (.ZN (n_3689), .A1 (inputA[15]), .A2 (inputB[25]));
NOR2_X1 i_4163 (.ZN (n_3687), .A1 (n_3697), .A2 (n_3689));
INV_X1 i_4162 (.ZN (n_3683), .A (n_3687));
AOI22_X1 i_4161 (.ZN (n_3682), .A1 (inputA[15]), .A2 (inputB[24]), .B1 (inputA[14]), .B2 (inputB[25]));
NOR2_X1 i_4160 (.ZN (n_3681), .A1 (n_3687), .A2 (n_3682));
NAND2_X1 i_4159 (.ZN (n_3680), .A1 (inputA[16]), .A2 (inputB[23]));
AOI21_X1 i_4158 (.ZN (n_3679), .A (n_3682), .B1 (n_3683), .B2 (n_3680));
OAI22_X1 i_4157 (.ZN (n_3678), .A1 (n_3718), .A2 (n_3717), .B1 (n_3716), .B2 (n_3715));
XOR2_X1 i_4156 (.Z (n_3677), .A (n_3679), .B (n_3678));
NAND2_X1 i_4155 (.ZN (n_3676), .A1 (inputA[12]), .A2 (inputB[26]));
NAND2_X1 i_4154 (.ZN (n_3675), .A1 (inputA[13]), .A2 (inputB[27]));
NOR2_X1 i_4153 (.ZN (n_3674), .A1 (n_3676), .A2 (n_3675));
AOI22_X1 i_4152 (.ZN (n_3673), .A1 (inputA[12]), .A2 (inputB[27]), .B1 (inputA[13]), .B2 (inputB[26]));
NOR2_X1 i_4151 (.ZN (n_3672), .A1 (n_3674), .A2 (n_3673));
NOR2_X1 i_4150 (.ZN (n_3671), .A1 (n_127), .A2 (n_1136));
AOI21_X1 i_4149 (.ZN (n_3670), .A (n_3674), .B1 (n_3672), .B2 (n_3671));
INV_X1 i_4148 (.ZN (n_3669), .A (n_3670));
AOI22_X1 i_4147 (.ZN (n_3642), .A1 (n_3679), .A2 (n_3678), .B1 (n_3677), .B2 (n_3669));
INV_X1 i_4146 (.ZN (n_3641), .A (n_3642));
XNOR2_X1 i_4145 (.ZN (n_3640), .A (n_3777), .B (n_3675));
NAND2_X1 i_4144 (.ZN (n_3639), .A1 (inputA[12]), .A2 (inputB[28]));
NAND2_X1 i_4143 (.ZN (n_3638), .A1 (inputA[11]), .A2 (inputB[29]));
AND2_X1 i_4142 (.ZN (n_3637), .A1 (inputA[9]), .A2 (inputB[31]));
XOR2_X1 i_4141 (.Z (n_3636), .A (n_3638), .B (n_3637));
INV_X1 i_4140 (.ZN (n_3632), .A (n_3636));
NAND2_X1 i_4139 (.ZN (n_3631), .A1 (inputA[10]), .A2 (inputB[30]));
OAI22_X1 i_4138 (.ZN (n_3630), .A1 (n_3777), .A2 (n_3675), .B1 (n_3640), .B2 (n_3639));
OAI22_X1 i_4137 (.ZN (n_3629), .A1 (n_3638), .A2 (n_3637), .B1 (n_3632), .B2 (n_3631));
XOR2_X1 i_4136 (.Z (n_3628), .A (n_3630), .B (n_3629));
AOI22_X1 i_4135 (.ZN (n_3627), .A1 (n_3630), .A2 (n_3629), .B1 (n_3641), .B2 (n_3628));
AOI21_X1 i_4134 (.ZN (n_3626), .A (n_3722), .B1 (n_3721), .B2 (n_3627));
NAND2_X1 i_4133 (.ZN (n_3625), .A1 (inputB[15]), .A2 (inputA[27]));
NAND2_X1 i_4132 (.ZN (n_3624), .A1 (inputB[14]), .A2 (inputA[28]));
XNOR2_X1 i_4131 (.ZN (n_3623), .A (n_3625), .B (n_3624));
NOR2_X1 i_4130 (.ZN (n_3622), .A1 (n_881), .A2 (n_585));
NAND3_X1 i_4129 (.ZN (n_3621), .A1 (inputB[18]), .A2 (n_3622), .A3 (inputA[25]));
INV_X1 i_4128 (.ZN (n_3620), .A (n_3621));
AOI22_X1 i_4127 (.ZN (n_3619), .A1 (inputB[18]), .A2 (inputA[24]), .B1 (inputB[17]), .B2 (inputA[25]));
NOR2_X1 i_4126 (.ZN (n_3618), .A1 (n_3620), .A2 (n_3619));
NAND2_X1 i_4125 (.ZN (n_3613), .A1 (inputB[19]), .A2 (inputA[23]));
OAI33_X1 i_4124 (.ZN (n_3612), .A1 (n_588), .A2 (n_214), .A3 (n_3623), .B1 (n_587)
    , .B2 (n_215), .B3 (n_3624));
OAI21_X1 i_4122 (.ZN (n_3611), .A (n_3621), .B1 (n_3619), .B2 (n_3613));
XOR2_X1 i_4121 (.Z (n_3610), .A (n_3612), .B (n_3611));
NAND2_X1 i_4120 (.ZN (n_3609), .A1 (inputB[21]), .A2 (inputA[21]));
NAND2_X1 i_4119 (.ZN (n_3608), .A1 (inputB[20]), .A2 (inputA[22]));
XNOR2_X1 i_4118 (.ZN (n_3607), .A (n_3609), .B (n_3608));
NAND2_X1 i_4117 (.ZN (n_3606), .A1 (inputB[22]), .A2 (inputA[20]));
OAI22_X1 i_4116 (.ZN (n_3605), .A1 (n_3609), .A2 (n_3608), .B1 (n_3607), .B2 (n_3606));
AOI22_X1 i_4115 (.ZN (n_3604), .A1 (n_3612), .A2 (n_3611), .B1 (n_3610), .B2 (n_3605));
NAND2_X1 i_4114 (.ZN (n_3603), .A1 (inputB[27]), .A2 (inputA[15]));
NAND2_X1 i_4113 (.ZN (n_3602), .A1 (inputB[26]), .A2 (inputA[16]));
XNOR2_X1 i_4112 (.ZN (n_3601), .A (n_3603), .B (n_3602));
NAND2_X1 i_4111 (.ZN (n_3598), .A1 (inputB[28]), .A2 (inputA[14]));
NAND2_X1 i_4110 (.ZN (n_3597), .A1 (inputB[24]), .A2 (inputA[17]));
NAND2_X1 i_4109 (.ZN (n_3596), .A1 (inputB[25]), .A2 (inputA[18]));
NOR2_X1 i_4108 (.ZN (n_3595), .A1 (n_3597), .A2 (n_3596));
AOI22_X1 i_4107 (.ZN (n_3594), .A1 (inputB[25]), .A2 (inputA[17]), .B1 (inputB[24]), .B2 (inputA[18]));
NOR2_X1 i_4106 (.ZN (n_3593), .A1 (n_3595), .A2 (n_3594));
NOR2_X1 i_4105 (.ZN (n_3592), .A1 (n_480), .A2 (n_218));
AOI21_X1 i_4104 (.ZN (n_3591), .A (n_3595), .B1 (n_3593), .B2 (n_3592));
INV_X1 i_4103 (.ZN (n_3590), .A (n_3591));
OAI22_X1 i_4102 (.ZN (n_3589), .A1 (n_3603), .A2 (n_3602), .B1 (n_3601), .B2 (n_3598));
XOR2_X1 i_4101 (.Z (n_3588), .A (n_3590), .B (n_3589));
NOR2_X1 i_4100 (.ZN (n_3587), .A1 (n_1136), .A2 (n_129));
NAND2_X1 i_4099 (.ZN (n_3586), .A1 (inputB[29]), .A2 (inputA[13]));
XNOR2_X1 i_4098 (.ZN (n_3585), .A (n_3587), .B (n_3586));
NAND2_X1 i_4097 (.ZN (n_3584), .A1 (inputB[30]), .A2 (inputA[12]));
OAI22_X1 i_4096 (.ZN (n_3572), .A1 (n_3587), .A2 (n_3586), .B1 (n_3585), .B2 (n_3584));
AOI22_X1 i_4095 (.ZN (n_3571), .A1 (n_3590), .A2 (n_3589), .B1 (n_3588), .B2 (n_3572));
NOR2_X1 i_4094 (.ZN (n_3570), .A1 (n_494), .A2 (n_3586));
AOI22_X1 i_4093 (.ZN (n_3569), .A1 (inputB[29]), .A2 (inputA[14]), .B1 (inputB[30]), .B2 (inputA[13]));
NOR2_X1 i_4092 (.ZN (n_3568), .A1 (n_3570), .A2 (n_3569));
NAND2_X1 i_4091 (.ZN (n_3567), .A1 (inputB[31]), .A2 (inputA[12]));
AOI21_X1 i_4090 (.ZN (n_3566), .A (n_3570), .B1 (n_3568), .B2 (n_3567));
XOR2_X1 i_4089 (.Z (n_3565), .A (n_3571), .B (n_3566));
XOR2_X1 i_4088 (.Z (n_3564), .A (n_3604), .B (n_3565));
NAND2_X1 i_4087 (.ZN (n_3563), .A1 (inputB[2]), .A2 (inputA[23]));
XNOR2_X1 i_4086 (.ZN (n_3562), .A (n_2969), .B (n_3563));
NOR2_X1 i_4085 (.ZN (n_3545), .A1 (n_2818), .A2 (n_2954));
AOI22_X1 i_4084 (.ZN (n_3544), .A1 (inputB[6]), .A2 (inputA[19]), .B1 (inputB[5]), .B2 (inputA[20]));
NOR2_X1 i_4083 (.ZN (n_3543), .A1 (n_3545), .A2 (n_3544));
OAI33_X1 i_4082 (.ZN (n_3542), .A1 (n_690), .A2 (n_482), .A3 (n_3562), .B1 (n_2925)
    , .B2 (n_685), .B3 (n_213));
OAI22_X1 i_4081 (.ZN (n_3541), .A1 (n_2818), .A2 (n_2954), .B1 (n_2959), .B2 (n_3544));
XOR2_X1 i_4080 (.Z (n_3540), .A (n_3542), .B (n_3541));
NAND2_X1 i_4079 (.ZN (n_3539), .A1 (inputB[10]), .A2 (inputA[15]));
XNOR2_X1 i_4078 (.ZN (n_3538), .A (n_2824), .B (n_3539));
NAND2_X1 i_4077 (.ZN (n_3537), .A1 (inputB[8]), .A2 (inputA[17]));
OAI22_X1 i_4076 (.ZN (n_3536), .A1 (n_2824), .A2 (n_3539), .B1 (n_3538), .B2 (n_3537));
AOI22_X1 i_4075 (.ZN (n_3535), .A1 (n_3542), .A2 (n_3541), .B1 (n_3540), .B2 (n_3536));
INV_X1 i_4074 (.ZN (n_3534), .A (n_2849));
NOR2_X1 i_4073 (.ZN (n_3525), .A1 (n_2848), .A2 (n_3043));
AOI22_X1 i_4072 (.ZN (n_3519), .A1 (inputA[6]), .A2 (inputB[19]), .B1 (inputA[7]), .B2 (inputB[18]));
NOR2_X1 i_4071 (.ZN (n_3518), .A1 (n_3525), .A2 (n_3519));
NAND2_X1 i_4070 (.ZN (n_3517), .A1 (n_3534), .A2 (n_3518));
AOI21_X1 i_4069 (.ZN (n_3516), .A (n_3525), .B1 (n_3534), .B2 (n_3518));
NOR3_X1 i_4068 (.ZN (n_3512), .A1 (n_2787), .A2 (n_530), .A3 (n_880));
AOI22_X1 i_4067 (.ZN (n_3511), .A1 (inputA[14]), .A2 (inputB[11]), .B1 (inputA[13]), .B2 (inputB[12]));
NOR2_X1 i_4066 (.ZN (n_3510), .A1 (n_3512), .A2 (n_3511));
NOR2_X1 i_4065 (.ZN (n_3509), .A1 (n_667), .A2 (n_671));
AOI21_X1 i_4064 (.ZN (n_3508), .A (n_3512), .B1 (n_3510), .B2 (n_3509));
XNOR2_X1 i_4063 (.ZN (n_3507), .A (n_3516), .B (n_3508));
XOR2_X1 i_4062 (.Z (n_3506), .A (n_3022), .B (n_3020));
XOR2_X1 i_4061 (.Z (n_3501), .A (n_3386), .B (n_3383));
XOR2_X1 i_4060 (.Z (n_3500), .A (n_3506), .B (n_3501));
XOR2_X1 i_4059 (.Z (n_3499), .A (n_3026), .B (n_3025));
AOI22_X1 i_4058 (.ZN (n_3498), .A1 (n_3506), .A2 (n_3501), .B1 (n_3500), .B2 (n_3499));
XNOR2_X1 i_4057 (.ZN (n_3497), .A (n_3371), .B (n_3360));
XOR2_X1 i_4056 (.Z (n_3496), .A (n_3498), .B (n_3497));
XOR2_X1 i_4055 (.Z (n_3493), .A (n_3370), .B (n_3361));
XNOR2_X1 i_4054 (.ZN (n_3492), .A (n_3397), .B (n_2944));
XOR2_X1 i_4053 (.Z (n_3491), .A (n_3493), .B (n_3492));
XNOR2_X1 i_4052 (.ZN (n_3490), .A (n_3399), .B (n_21));
NAND2_X1 i_4051 (.ZN (n_3489), .A1 (n_3491), .A2 (n_3490));
OAI21_X1 i_4049 (.ZN (n_3488), .A (n_3489), .B1 (n_3493), .B2 (n_3492));
AOI22_X1 i_4048 (.ZN (n_3487), .A1 (n_3498), .A2 (n_3497), .B1 (n_3496), .B2 (n_3488));
XNOR2_X1 i_4047 (.ZN (n_3486), .A (n_3356), .B (n_3355));
XOR2_X1 i_4046 (.Z (n_3485), .A (n_3487), .B (n_3486));
OAI22_X1 i_4045 (.ZN (n_3484), .A1 (n_3507), .A2 (n_17), .B1 (n_3516), .B2 (n_3508));
OAI22_X1 i_4044 (.ZN (n_3483), .A1 (n_2708), .A2 (n_2707), .B1 (n_2711), .B2 (n_2710));
NOR2_X1 i_4043 (.ZN (n_3482), .A1 (n_3484), .A2 (n_3483));
AOI21_X1 i_4042 (.ZN (n_3481), .A (n_3482), .B1 (n_3484), .B2 (n_3483));
INV_X1 i_4041 (.ZN (n_3480), .A (n_3481));
AOI21_X1 i_4040 (.ZN (n_3479), .A (n_3482), .B1 (n_3535), .B2 (n_3481));
XOR2_X1 i_4039 (.Z (n_3478), .A (n_3031), .B (n_3017));
XNOR2_X1 i_4038 (.ZN (n_3477), .A (n_3479), .B (n_3478));
XOR2_X1 i_4037 (.Z (n_3476), .A (n_3392), .B (n_3382));
INV_X1 i_4036 (.ZN (n_3475), .A (n_3476));
OAI22_X1 i_4035 (.ZN (n_3474), .A1 (n_3479), .A2 (n_3478), .B1 (n_3477), .B2 (n_3476));
INV_X1 i_4034 (.ZN (n_3473), .A (n_3474));
AOI22_X1 i_4033 (.ZN (n_3472), .A1 (n_3487), .A2 (n_3486), .B1 (n_3485), .B2 (n_3473));
XNOR2_X1 i_4032 (.ZN (n_3471), .A (n_3423), .B (n_3416));
NOR2_X1 i_4031 (.ZN (n_3470), .A1 (n_3472), .A2 (n_3471));
AOI21_X1 i_4030 (.ZN (n_3469), .A (n_3470), .B1 (n_3472), .B2 (n_3471));
OAI21_X1 i_4029 (.ZN (n_3468), .A (n_3237), .B1 (n_3285), .B2 (n_3238));
AOI21_X1 i_4028 (.ZN (n_3467), .A (n_3470), .B1 (n_3469), .B2 (n_3468));
XOR2_X1 i_4027 (.Z (n_3466), .A (n_1698), .B (n_1697));
XOR2_X1 i_4026 (.Z (n_3465), .A (n_1704), .B (n_1703));
XOR2_X1 i_4025 (.Z (n_3464), .A (n_3466), .B (n_3465));
XOR2_X1 i_4024 (.Z (n_3463), .A (n_1680), .B (n_1679));
AOI22_X1 i_4023 (.ZN (n_3462), .A1 (n_3466), .A2 (n_3465), .B1 (n_3464), .B2 (n_3463));
XOR2_X1 i_4022 (.Z (n_3461), .A (n_3428), .B (n_3414));
NOR2_X1 i_4021 (.ZN (n_3460), .A1 (n_3462), .A2 (n_3461));
AOI21_X1 i_4020 (.ZN (n_3459), .A (n_3460), .B1 (n_3462), .B2 (n_3461));
AOI21_X1 i_4019 (.ZN (n_3458), .A (n_3460), .B1 (n_3467), .B2 (n_3459));
XNOR2_X1 i_4018 (.ZN (n_3457), .A (n_3324), .B (n_3296));
NOR2_X1 i_4017 (.ZN (n_3456), .A1 (n_3458), .A2 (n_3457));
AOI21_X1 i_4016 (.ZN (n_3455), .A (n_3456), .B1 (n_3458), .B2 (n_3457));
XNOR2_X1 i_4015 (.ZN (n_3454), .A (n_3410), .B (n_3409));
AOI21_X1 i_4014 (.ZN (n_3453), .A (n_3456), .B1 (n_3455), .B2 (n_3454));
INV_X1 i_4013 (.ZN (n_3452), .A (n_3286));
INV_X1 i_4012 (.ZN (n_3451), .A (n_2953));
INV_X1 i_4011 (.ZN (n_3433), .A (n_3172));
INV_X1 i_4010 (.ZN (n_3432), .A (n_2929));
INV_X1 i_4009 (.ZN (n_3431), .A (n_2937));
OAI21_X1 i_4008 (.ZN (n_3430), .A (n_3288), .B1 (n_3452), .B2 (n_3287));
XOR2_X1 i_4007 (.Z (n_3429), .A (n_1294), .B (n_1285));
XOR2_X1 i_4006 (.Z (n_3428), .A (n_3430), .B (n_3429));
XOR2_X1 i_4005 (.Z (n_3426), .A (n_1289), .B (n_1286));
XOR2_X1 i_4004 (.Z (n_3425), .A (n_1309), .B (n_1308));
NOR2_X1 i_4003 (.ZN (n_3424), .A1 (n_3426), .A2 (n_3425));
AOI21_X1 i_4002 (.ZN (n_3423), .A (n_3424), .B1 (n_3426), .B2 (n_3425));
XOR2_X1 i_4001 (.Z (n_3422), .A (n_29), .B (n_30));
XOR2_X1 i_4000 (.Z (n_3421), .A (n_1302), .B (n_1301));
NOR2_X1 i_3999 (.ZN (n_3420), .A1 (n_3422), .A2 (n_3421));
AOI21_X1 i_3998 (.ZN (n_3418), .A (n_3420), .B1 (n_3422), .B2 (n_3421));
XNOR2_X1 i_3997 (.ZN (n_3417), .A (n_1595), .B (n_1594));
AOI21_X1 i_3996 (.ZN (n_3416), .A (n_3420), .B1 (n_3418), .B2 (n_3417));
INV_X1 i_3995 (.ZN (n_3415), .A (n_3416));
AOI21_X1 i_3994 (.ZN (n_3414), .A (n_3424), .B1 (n_3423), .B2 (n_3415));
INV_X1 i_3993 (.ZN (n_3413), .A (n_3414));
AOI22_X1 i_3992 (.ZN (n_3412), .A1 (n_3430), .A2 (n_3429), .B1 (n_3428), .B2 (n_3413));
XOR2_X1 i_3991 (.Z (n_3411), .A (n_1240), .B (n_1229));
XOR2_X1 i_3990 (.Z (n_3410), .A (n_3412), .B (n_3411));
XOR2_X1 i_3989 (.Z (n_3409), .A (n_1282), .B (n_1281));
AOI22_X1 i_3988 (.ZN (n_3408), .A1 (n_3412), .A2 (n_3411), .B1 (n_3410), .B2 (n_3409));
XNOR2_X1 i_3987 (.ZN (n_3407), .A (n_1226), .B (n_1280));
XNOR2_X1 i_3986 (.ZN (n_3400), .A (n_3408), .B (n_3407));
XNOR2_X1 i_3985 (.ZN (n_3399), .A (n_3051), .B (n_20));
NOR2_X1 i_3984 (.ZN (n_3398), .A1 (n_2940), .A2 (n_3178));
NOR2_X1 i_3983 (.ZN (n_3397), .A1 (n_19), .A2 (n_3398));
OAI33_X1 i_3982 (.ZN (n_3394), .A1 (n_1894), .A2 (n_400), .A3 (n_3399), .B1 (n_3051)
    , .B2 (n_1136), .B3 (n_588));
OAI22_X1 i_3981 (.ZN (n_3393), .A1 (n_2940), .A2 (n_3178), .B1 (n_19), .B2 (n_2944));
XOR2_X1 i_3980 (.Z (n_3392), .A (n_3394), .B (n_3393));
NOR2_X1 i_3979 (.ZN (n_3391), .A1 (n_864), .A2 (n_414));
NOR2_X1 i_3978 (.ZN (n_3390), .A1 (n_1551), .A2 (n_314));
NAND2_X1 i_3977 (.ZN (n_3387), .A1 (n_3391), .A2 (n_3390));
OAI21_X1 i_3976 (.ZN (n_3386), .A (n_3387), .B1 (n_3391), .B2 (n_3390));
NAND2_X1 i_3975 (.ZN (n_3383), .A1 (inputA[6]), .A2 (inputB[21]));
OAI21_X1 i_3974 (.ZN (n_3382), .A (n_3387), .B1 (n_3386), .B2 (n_3383));
NOR2_X1 i_3973 (.ZN (n_3381), .A1 (n_2963), .A2 (n_3148));
NAND2_X1 i_3972 (.ZN (n_3378), .A1 (inputA[20]), .A2 (inputB[7]));
XNOR2_X1 i_3971 (.ZN (n_3377), .A (n_2958), .B (n_3378));
NAND2_X1 i_3970 (.ZN (n_3376), .A1 (inputA[18]), .A2 (inputB[9]));
OAI21_X1 i_3969 (.ZN (n_3374), .A (n_18), .B1 (n_2963), .B2 (n_3148));
OAI22_X1 i_3968 (.ZN (n_3373), .A1 (n_2958), .A2 (n_3378), .B1 (n_3377), .B2 (n_3376));
NAND2_X1 i_3966 (.ZN (n_3372), .A1 (n_3374), .A2 (n_3373));
OAI21_X1 i_3965 (.ZN (n_3371), .A (n_3372), .B1 (n_3374), .B2 (n_3373));
AOI22_X1 i_3964 (.ZN (n_3370), .A1 (n_3451), .A2 (n_3433), .B1 (n_2953), .B2 (n_3172));
NOR2_X1 i_3963 (.ZN (n_3361), .A1 (n_880), .A2 (n_478));
AOI22_X1 i_3962 (.ZN (n_3360), .A1 (n_3451), .A2 (n_3433), .B1 (n_3370), .B2 (n_3361));
AOI22_X1 i_3961 (.ZN (n_3359), .A1 (n_3394), .A2 (n_3393), .B1 (n_3392), .B2 (n_3382));
INV_X1 i_3960 (.ZN (n_3358), .A (n_3359));
OAI21_X1 i_3959 (.ZN (n_3357), .A (n_3372), .B1 (n_3371), .B2 (n_3360));
XOR2_X1 i_3958 (.Z (n_3356), .A (n_3358), .B (n_3357));
AOI22_X1 i_3957 (.ZN (n_3355), .A1 (n_2932), .A2 (n_2931), .B1 (n_3432), .B2 (n_2930));
INV_X1 i_3956 (.ZN (n_3354), .A (n_3355));
AOI22_X1 i_3955 (.ZN (n_3353), .A1 (n_3358), .A2 (n_3357), .B1 (n_3356), .B2 (n_3354));
XOR2_X1 i_3954 (.Z (n_3352), .A (n_1606), .B (n_1591));
XOR2_X1 i_3953 (.Z (n_3351), .A (n_1304), .B (n_1300));
NOR2_X1 i_3952 (.ZN (n_3350), .A1 (n_3352), .A2 (n_3351));
AOI21_X1 i_3951 (.ZN (n_3349), .A (n_3350), .B1 (n_3352), .B2 (n_3351));
AOI21_X1 i_3950 (.ZN (n_3348), .A (n_3350), .B1 (n_3353), .B2 (n_3349));
XOR2_X1 i_3949 (.Z (n_3347), .A (n_1586), .B (n_1573));
XNOR2_X1 i_3948 (.ZN (n_3346), .A (n_1251), .B (n_1244));
XNOR2_X1 i_3947 (.ZN (n_3327), .A (n_3347), .B (n_3346));
OAI22_X1 i_3946 (.ZN (n_3326), .A1 (n_3347), .A2 (n_3346), .B1 (n_3348), .B2 (n_3327));
XNOR2_X1 i_3945 (.ZN (n_3325), .A (n_1648), .B (n_1563));
XOR2_X1 i_3944 (.Z (n_3324), .A (n_3326), .B (n_3325));
AOI22_X1 i_3943 (.ZN (n_3323), .A1 (n_3013), .A2 (n_3012), .B1 (n_3011), .B2 (n_3009));
AOI22_X1 i_3942 (.ZN (n_3320), .A1 (n_3431), .A2 (n_2960), .B1 (n_2936), .B2 (n_2928));
XOR2_X1 i_3941 (.Z (n_3319), .A (n_3134), .B (n_3133));
XNOR2_X1 i_3940 (.ZN (n_3318), .A (n_3104), .B (n_3103));
XOR2_X1 i_3939 (.Z (n_3316), .A (n_3319), .B (n_3318));
XNOR2_X1 i_3938 (.ZN (n_3315), .A (n_3146), .B (n_3145));
AOI22_X1 i_3937 (.ZN (n_3314), .A1 (n_3194), .A2 (n_3193), .B1 (n_3184), .B2 (n_3183));
AOI22_X1 i_3936 (.ZN (n_3313), .A1 (n_3319), .A2 (n_3318), .B1 (n_3316), .B2 (n_3315));
XNOR2_X1 i_3935 (.ZN (n_3312), .A (n_3314), .B (n_3313));
AOI22_X1 i_3934 (.ZN (n_3303), .A1 (n_3149), .A2 (n_3099), .B1 (n_3098), .B2 (n_3073));
OAI22_X1 i_3933 (.ZN (n_3302), .A1 (n_3314), .A2 (n_3313), .B1 (n_3320), .B2 (n_3312));
XOR2_X1 i_3932 (.Z (n_3301), .A (n_3303), .B (n_3302));
AOI22_X1 i_3931 (.ZN (n_3300), .A1 (n_3303), .A2 (n_3302), .B1 (n_3323), .B2 (n_3301));
XNOR2_X1 i_3930 (.ZN (n_3299), .A (n_1231), .B (n_1230));
XOR2_X1 i_3929 (.Z (n_3298), .A (n_1569), .B (n_1568));
XOR2_X1 i_3928 (.Z (n_3297), .A (n_3299), .B (n_3298));
AOI22_X1 i_3927 (.ZN (n_3296), .A1 (n_3299), .A2 (n_3298), .B1 (n_3300), .B2 (n_3297));
AOI22_X1 i_3926 (.ZN (n_3295), .A1 (n_3326), .A2 (n_3325), .B1 (n_3324), .B2 (n_3296));
XOR2_X1 i_3925 (.Z (n_3294), .A (n_3400), .B (n_3295));
INV_X1 i_3924 (.ZN (n_3293), .A (n_3151));
INV_X1 i_3923 (.ZN (n_3292), .A (n_3102));
XNOR2_X1 i_3922 (.ZN (n_3291), .A (n_1708), .B (n_1707));
AOI22_X1 i_3921 (.ZN (n_3290), .A1 (n_3293), .A2 (n_3156), .B1 (n_3174), .B2 (n_3157));
XNOR2_X1 i_3920 (.ZN (n_3289), .A (n_1334), .B (n_1333));
NAND2_X1 i_3919 (.ZN (n_3288), .A1 (n_3290), .A2 (n_3289));
OAI21_X1 i_3918 (.ZN (n_3287), .A (n_3288), .B1 (n_3290), .B2 (n_3289));
AOI22_X1 i_3917 (.ZN (n_3286), .A1 (n_3292), .A2 (n_3131), .B1 (n_3144), .B2 (n_3132));
XNOR2_X1 i_3916 (.ZN (n_3285), .A (n_3287), .B (n_3286));
NOR2_X1 i_3915 (.ZN (n_3284), .A1 (n_2929), .A2 (n_1340));
AOI22_X1 i_3914 (.ZN (n_3283), .A1 (inputB[1]), .A2 (inputA[28]), .B1 (inputB[0]), .B2 (inputA[29]));
NOR2_X1 i_3913 (.ZN (n_3281), .A1 (n_3284), .A2 (n_3283));
NOR2_X1 i_3912 (.ZN (n_3280), .A1 (n_1219), .A2 (n_215));
NOR2_X1 i_3911 (.ZN (n_3279), .A1 (n_3133), .A2 (n_1214));
AOI22_X1 i_3910 (.ZN (n_3278), .A1 (inputB[4]), .A2 (inputA[25]), .B1 (inputB[5]), .B2 (inputA[24]));
NOR2_X1 i_3909 (.ZN (n_3277), .A1 (n_3279), .A2 (n_3278));
XOR2_X1 i_3908 (.Z (n_3276), .A (n_3281), .B (n_3280));
XNOR2_X1 i_3907 (.ZN (n_3275), .A (n_3138), .B (n_3277));
NOR2_X1 i_3906 (.ZN (n_3274), .A1 (n_3276), .A2 (n_3275));
AOI21_X1 i_3905 (.ZN (n_3273), .A (n_3274), .B1 (n_3276), .B2 (n_3275));
NOR2_X1 i_3904 (.ZN (n_3272), .A1 (n_3148), .A2 (n_1441));
AOI22_X1 i_3903 (.ZN (n_3271), .A1 (inputB[7]), .A2 (inputA[22]), .B1 (inputB[6]), .B2 (inputA[23]));
NOR2_X1 i_3902 (.ZN (n_3270), .A1 (n_3272), .A2 (n_3271));
NOR2_X1 i_3901 (.ZN (n_3269), .A1 (n_669), .A2 (n_482));
XNOR2_X1 i_3900 (.ZN (n_3268), .A (n_3270), .B (n_3269));
NAND2_X1 i_3899 (.ZN (n_3256), .A1 (n_3273), .A2 (n_3268));
XNOR2_X1 i_3898 (.ZN (n_3255), .A (n_3107), .B (n_1432));
NAND2_X1 i_3897 (.ZN (n_3254), .A1 (inputB[11]), .A2 (inputA[18]));
NOR2_X1 i_3896 (.ZN (n_3253), .A1 (n_3178), .A2 (n_1472));
AOI22_X1 i_3895 (.ZN (n_3252), .A1 (inputB[16]), .A2 (inputA[13]), .B1 (inputB[15]), .B2 (inputA[14]));
NOR2_X1 i_3894 (.ZN (n_3251), .A1 (n_3253), .A2 (n_3252));
NAND2_X1 i_3893 (.ZN (n_3250), .A1 (n_1487), .A2 (n_3251));
OAI21_X1 i_3892 (.ZN (n_3249), .A (n_3250), .B1 (n_1487), .B2 (n_3251));
XNOR2_X1 i_3891 (.ZN (n_3248), .A (n_3255), .B (n_3254));
XOR2_X1 i_3890 (.Z (n_3247), .A (n_3249), .B (n_3248));
XNOR2_X1 i_3889 (.ZN (n_3246), .A (n_1288), .B (n_1287));
AOI21_X1 i_3888 (.ZN (n_3245), .A (n_3274), .B1 (n_3273), .B2 (n_3268));
AOI22_X1 i_3885 (.ZN (n_3244), .A1 (n_3249), .A2 (n_3248), .B1 (n_3247), .B2 (n_3246));
XOR2_X1 i_3884 (.Z (n_3238), .A (n_3245), .B (n_3244));
NAND2_X1 i_3883 (.ZN (n_3237), .A1 (n_3285), .A2 (n_3238));
OAI21_X1 i_3882 (.ZN (n_3236), .A (n_3237), .B1 (n_3245), .B2 (n_3244));
XOR2_X1 i_3881 (.Z (n_3235), .A (n_3291), .B (n_3236));
XNOR2_X1 i_3880 (.ZN (n_3234), .A (n_1689), .B (n_1678));
XNOR2_X1 i_3879 (.ZN (n_3233), .A (n_3235), .B (n_3234));
INV_X1 i_3878 (.ZN (n_3232), .A (n_2834));
OAI21_X1 i_3877 (.ZN (n_3218), .A (n_2839), .B1 (n_3232), .B2 (n_2838));
NOR2_X1 i_3876 (.ZN (n_3217), .A1 (n_2837), .A2 (n_2705));
AOI22_X1 i_3875 (.ZN (n_3216), .A1 (inputA[5]), .A2 (inputB[20]), .B1 (inputA[4]), .B2 (inputB[21]));
NOR2_X1 i_3874 (.ZN (n_3215), .A1 (n_3217), .A2 (n_3216));
NOR2_X1 i_3873 (.ZN (n_3214), .A1 (n_1724), .A2 (n_217));
OAI22_X1 i_3872 (.ZN (n_3213), .A1 (n_2829), .A2 (n_2828), .B1 (n_2763), .B2 (n_2830));
INV_X1 i_3871 (.ZN (n_3209), .A (n_3213));
AOI21_X1 i_3870 (.ZN (n_3208), .A (n_3217), .B1 (n_3215), .B2 (n_3214));
NOR2_X1 i_3869 (.ZN (n_3207), .A1 (n_3209), .A2 (n_3208));
AOI21_X1 i_3868 (.ZN (n_3206), .A (n_3207), .B1 (n_3209), .B2 (n_3208));
AOI21_X1 i_3867 (.ZN (n_3205), .A (n_3207), .B1 (n_3218), .B2 (n_3206));
XNOR2_X1 i_3866 (.ZN (n_3204), .A (n_3033), .B (n_3032));
NOR2_X1 i_3865 (.ZN (n_3201), .A1 (n_3205), .A2 (n_3204));
AOI21_X1 i_3864 (.ZN (n_3200), .A (n_3201), .B1 (n_3205), .B2 (n_3204));
XOR2_X1 i_3863 (.Z (n_3199), .A (n_2945), .B (n_2938));
AOI21_X1 i_3862 (.ZN (n_3198), .A (n_3201), .B1 (n_3200), .B2 (n_3199));
XOR2_X1 i_3861 (.Z (n_3196), .A (n_3074), .B (n_3075));
XOR2_X1 i_3860 (.Z (n_3195), .A (n_3198), .B (n_3196));
XOR2_X1 i_3859 (.Z (n_3194), .A (n_3169), .B (n_3168));
XNOR2_X1 i_3858 (.ZN (n_3193), .A (n_3176), .B (n_3175));
XOR2_X1 i_3857 (.Z (n_3184), .A (n_3194), .B (n_3193));
XNOR2_X1 i_3856 (.ZN (n_3183), .A (n_3153), .B (n_3152));
XOR2_X1 i_3855 (.Z (n_3182), .A (n_3184), .B (n_3183));
AOI22_X1 i_3854 (.ZN (n_3179), .A1 (n_3198), .A2 (n_3196), .B1 (n_3195), .B2 (n_3182));
NAND2_X1 i_3853 (.ZN (n_3178), .A1 (inputA[13]), .A2 (inputB[15]));
NAND2_X1 i_3852 (.ZN (n_3177), .A1 (inputA[14]), .A2 (inputB[14]));
XNOR2_X1 i_3851 (.ZN (n_3176), .A (n_3178), .B (n_3177));
NAND2_X1 i_3850 (.ZN (n_3175), .A1 (inputA[12]), .A2 (inputB[16]));
OAI22_X1 i_3849 (.ZN (n_3174), .A1 (n_3178), .A2 (n_3177), .B1 (n_3176), .B2 (n_3175));
NAND2_X1 i_3848 (.ZN (n_3172), .A1 (inputA[16]), .A2 (inputB[11]));
NOR2_X1 i_3847 (.ZN (n_3171), .A1 (n_1287), .A2 (n_3172));
AOI22_X1 i_3846 (.ZN (n_3170), .A1 (inputA[16]), .A2 (inputB[12]), .B1 (inputA[17]), .B2 (inputB[11]));
NOR2_X1 i_3845 (.ZN (n_3169), .A1 (n_3171), .A2 (n_3170));
NAND2_X1 i_3844 (.ZN (n_3168), .A1 (inputA[15]), .A2 (inputB[13]));
OAI22_X1 i_3843 (.ZN (n_3157), .A1 (n_1287), .A2 (n_3172), .B1 (n_3170), .B2 (n_3168));
XOR2_X1 i_3842 (.Z (n_3156), .A (n_3174), .B (n_3157));
NOR3_X1 i_3841 (.ZN (n_3155), .A1 (n_3051), .A2 (n_400), .A3 (n_1136));
AOI22_X1 i_3840 (.ZN (n_3154), .A1 (inputA[10]), .A2 (inputB[18]), .B1 (inputA[11]), .B2 (inputB[17]));
NOR2_X1 i_3839 (.ZN (n_3153), .A1 (n_3155), .A2 (n_3154));
NOR2_X1 i_3838 (.ZN (n_3152), .A1 (n_1894), .A2 (n_314));
AOI21_X1 i_3837 (.ZN (n_3151), .A (n_3155), .B1 (n_3153), .B2 (n_3152));
XOR2_X1 i_3836 (.Z (n_3150), .A (n_3156), .B (n_3151));
INV_X1 i_3835 (.ZN (n_3149), .A (n_3150));
NAND2_X1 i_3834 (.ZN (n_3148), .A1 (inputA[22]), .A2 (inputB[6]));
NAND2_X1 i_3833 (.ZN (n_3147), .A1 (inputA[21]), .A2 (inputB[7]));
XNOR2_X1 i_3832 (.ZN (n_3146), .A (n_3148), .B (n_3147));
NAND2_X1 i_3831 (.ZN (n_3145), .A1 (inputA[23]), .A2 (inputB[5]));
OAI22_X1 i_3830 (.ZN (n_3144), .A1 (n_3148), .A2 (n_3147), .B1 (n_3146), .B2 (n_3145));
NAND2_X1 i_3829 (.ZN (n_3138), .A1 (inputA[26]), .A2 (inputB[3]));
NOR2_X1 i_3828 (.ZN (n_3137), .A1 (n_2935), .A2 (n_3138));
AOI22_X1 i_3827 (.ZN (n_3136), .A1 (inputA[26]), .A2 (inputB[2]), .B1 (inputA[25]), .B2 (inputB[3]));
NOR2_X1 i_3826 (.ZN (n_3134), .A1 (n_3137), .A2 (n_3136));
NAND2_X1 i_3825 (.ZN (n_3133), .A1 (inputA[24]), .A2 (inputB[4]));
OAI22_X1 i_3824 (.ZN (n_3132), .A1 (n_2935), .A2 (n_3138), .B1 (n_3136), .B2 (n_3133));
XOR2_X1 i_3823 (.Z (n_3131), .A (n_3144), .B (n_3132));
NAND2_X1 i_3822 (.ZN (n_3107), .A1 (inputA[20]), .A2 (inputB[9]));
NOR2_X1 i_3821 (.ZN (n_3106), .A1 (n_2958), .A2 (n_3107));
AOI22_X1 i_3820 (.ZN (n_3105), .A1 (inputA[19]), .A2 (inputB[9]), .B1 (inputA[20]), .B2 (inputB[8]));
NOR2_X1 i_3819 (.ZN (n_3104), .A1 (n_3106), .A2 (n_3105));
NOR2_X1 i_3818 (.ZN (n_3103), .A1 (n_1131), .A2 (n_479));
AOI21_X1 i_3817 (.ZN (n_3102), .A (n_3106), .B1 (n_3104), .B2 (n_3103));
XOR2_X1 i_3816 (.Z (n_3101), .A (n_3131), .B (n_3102));
INV_X1 i_3815 (.ZN (n_3099), .A (n_3101));
AOI22_X1 i_3814 (.ZN (n_3098), .A1 (n_3150), .A2 (n_3101), .B1 (n_3149), .B2 (n_3099));
NAND2_X1 i_3813 (.ZN (n_3097), .A1 (inputA[6]), .A2 (inputB[22]));
XOR2_X1 i_3812 (.Z (n_3096), .A (n_1642), .B (n_3097));
XNOR2_X1 i_3811 (.ZN (n_3095), .A (n_1645), .B (n_1644));
XOR2_X1 i_3810 (.Z (n_3075), .A (n_3096), .B (n_3095));
XNOR2_X1 i_3809 (.ZN (n_3074), .A (n_1634), .B (n_1633));
AOI22_X1 i_3808 (.ZN (n_3073), .A1 (n_3096), .A2 (n_3095), .B1 (n_3075), .B2 (n_3074));
XNOR2_X1 i_3807 (.ZN (n_3072), .A (n_3098), .B (n_3073));
NAND2_X1 i_3806 (.ZN (n_3071), .A1 (inputA[9]), .A2 (inputB[16]));
NAND2_X1 i_3805 (.ZN (n_3051), .A1 (inputA[10]), .A2 (inputB[17]));
AOI22_X1 i_3804 (.ZN (n_3050), .A1 (inputA[10]), .A2 (inputB[16]), .B1 (inputA[9]), .B2 (inputB[17]));
INV_X1 i_3803 (.ZN (n_3049), .A (n_3050));
OAI21_X1 i_3801 (.ZN (n_3048), .A (n_3049), .B1 (n_3071), .B2 (n_3051));
NAND2_X1 i_3799 (.ZN (n_3047), .A1 (inputA[11]), .A2 (inputB[15]));
NAND2_X1 i_3798 (.ZN (n_3043), .A1 (inputA[7]), .A2 (inputB[19]));
NAND2_X1 i_3797 (.ZN (n_3042), .A1 (inputA[8]), .A2 (inputB[18]));
XNOR2_X1 i_3796 (.ZN (n_3040), .A (n_3043), .B (n_3042));
OAI33_X1 i_3795 (.ZN (n_3039), .A1 (n_1349), .A2 (n_414), .A3 (n_3040), .B1 (n_1551)
    , .B2 (n_400), .B3 (n_3043));
OAI22_X1 i_3794 (.ZN (n_3038), .A1 (n_3071), .A2 (n_3051), .B1 (n_3048), .B2 (n_3047));
XOR2_X1 i_3793 (.Z (n_3033), .A (n_3039), .B (n_3038));
OAI22_X1 i_3792 (.ZN (n_3032), .A1 (n_2702), .A2 (n_2701), .B1 (n_2705), .B2 (n_2704));
AOI22_X1 i_3791 (.ZN (n_3031), .A1 (n_3039), .A2 (n_3038), .B1 (n_3033), .B2 (n_3032));
NOR2_X1 i_3790 (.ZN (n_3030), .A1 (n_2711), .A2 (n_1638));
AOI22_X1 i_3789 (.ZN (n_3029), .A1 (inputA[1]), .A2 (inputB[26]), .B1 (inputA[2]), .B2 (inputB[25]));
NOR2_X1 i_3788 (.ZN (n_3026), .A1 (n_3030), .A2 (n_3029));
NOR2_X1 i_3787 (.ZN (n_3025), .A1 (n_66), .A2 (n_126));
NOR2_X1 i_3786 (.ZN (n_3024), .A1 (n_2704), .A2 (n_1647));
AOI22_X1 i_3785 (.ZN (n_3023), .A1 (inputA[4]), .A2 (inputB[23]), .B1 (inputA[5]), .B2 (inputB[22]));
NOR2_X1 i_3784 (.ZN (n_3022), .A1 (n_3024), .A2 (n_3023));
NOR2_X1 i_3783 (.ZN (n_3020), .A1 (n_1724), .A2 (n_461));
AOI21_X1 i_3782 (.ZN (n_3019), .A (n_3030), .B1 (n_3026), .B2 (n_3025));
AOI21_X1 i_3781 (.ZN (n_3018), .A (n_3024), .B1 (n_3022), .B2 (n_3020));
XNOR2_X1 i_3780 (.ZN (n_3017), .A (n_3019), .B (n_3018));
OAI22_X1 i_3779 (.ZN (n_3013), .A1 (n_3019), .A2 (n_3018), .B1 (n_3031), .B2 (n_3017));
XNOR2_X1 i_3778 (.ZN (n_3012), .A (n_1603), .B (n_1599));
XOR2_X1 i_3777 (.Z (n_3011), .A (n_3013), .B (n_3012));
XOR2_X1 i_3776 (.Z (n_3009), .A (n_1639), .B (n_1607));
XNOR2_X1 i_3775 (.ZN (n_3008), .A (n_3011), .B (n_3009));
NAND2_X1 i_3774 (.ZN (n_3007), .A1 (inputB[0]), .A2 (inputA[25]));
NAND2_X1 i_3773 (.ZN (n_2998), .A1 (inputB[1]), .A2 (inputA[26]));
NOR2_X1 i_3772 (.ZN (n_2990), .A1 (n_3007), .A2 (n_2998));
AOI22_X1 i_3771 (.ZN (n_2980), .A1 (inputB[1]), .A2 (inputA[25]), .B1 (inputB[0]), .B2 (inputA[26]));
NOR2_X1 i_3770 (.ZN (n_2979), .A1 (n_2990), .A2 (n_2980));
NOR2_X1 i_3769 (.ZN (n_2978), .A1 (n_1219), .A2 (n_585));
AOI21_X1 i_3768 (.ZN (n_2977), .A (n_2990), .B1 (n_2979), .B2 (n_2978));
NOR3_X1 i_3767 (.ZN (n_2976), .A1 (n_62), .A2 (n_215), .A3 (n_2977));
OAI21_X1 i_3766 (.ZN (n_2975), .A (n_2977), .B1 (n_62), .B2 (n_215));
INV_X1 i_3765 (.ZN (n_2971), .A (n_2975));
NOR2_X1 i_3764 (.ZN (n_2970), .A1 (n_2976), .A2 (n_2971));
NAND2_X1 i_3763 (.ZN (n_2969), .A1 (inputB[3]), .A2 (inputA[22]));
NAND2_X1 i_3762 (.ZN (n_2968), .A1 (inputB[4]), .A2 (inputA[23]));
NOR2_X1 i_3761 (.ZN (n_2967), .A1 (n_2969), .A2 (n_2968));
INV_X1 i_3760 (.ZN (n_2966), .A (n_2967));
AOI22_X1 i_3759 (.ZN (n_2965), .A1 (inputB[4]), .A2 (inputA[22]), .B1 (inputB[3]), .B2 (inputA[23]));
NOR2_X1 i_3758 (.ZN (n_2964), .A1 (n_2967), .A2 (n_2965));
NAND2_X1 i_3757 (.ZN (n_2963), .A1 (inputB[5]), .A2 (inputA[21]));
AOI21_X1 i_3756 (.ZN (n_2962), .A (n_2965), .B1 (n_2966), .B2 (n_2963));
INV_X1 i_3755 (.ZN (n_2961), .A (n_2962));
OAI21_X1 i_3754 (.ZN (n_2960), .A (n_2975), .B1 (n_2976), .B2 (n_2962));
NAND2_X1 i_3753 (.ZN (n_2959), .A1 (inputB[7]), .A2 (inputA[18]));
NAND2_X1 i_3752 (.ZN (n_2958), .A1 (inputB[8]), .A2 (inputA[19]));
AOI22_X1 i_3751 (.ZN (n_2957), .A1 (inputB[7]), .A2 (inputA[19]), .B1 (inputB[8]), .B2 (inputA[18]));
INV_X1 i_3750 (.ZN (n_2956), .A (n_2957));
OAI21_X1 i_3749 (.ZN (n_2955), .A (n_2956), .B1 (n_2959), .B2 (n_2958));
NAND2_X1 i_3748 (.ZN (n_2954), .A1 (inputB[6]), .A2 (inputA[20]));
NAND2_X1 i_3747 (.ZN (n_2953), .A1 (inputB[10]), .A2 (inputA[17]));
AOI22_X1 i_3746 (.ZN (n_2952), .A1 (inputB[10]), .A2 (inputA[16]), .B1 (inputB[9]), .B2 (inputA[17]));
INV_X1 i_3745 (.ZN (n_2951), .A (n_2952));
OAI21_X1 i_3744 (.ZN (n_2950), .A (n_2951), .B1 (n_2824), .B2 (n_2953));
NAND2_X1 i_3743 (.ZN (n_2949), .A1 (inputB[11]), .A2 (inputA[15]));
OAI22_X1 i_3742 (.ZN (n_2948), .A1 (n_2824), .A2 (n_2953), .B1 (n_2950), .B2 (n_2949));
OAI22_X1 i_3741 (.ZN (n_2947), .A1 (n_2959), .A2 (n_2958), .B1 (n_2955), .B2 (n_2954));
NAND2_X1 i_3740 (.ZN (n_2946), .A1 (n_2948), .A2 (n_2947));
OAI21_X1 i_3739 (.ZN (n_2945), .A (n_2946), .B1 (n_2948), .B2 (n_2947));
NAND2_X1 i_3738 (.ZN (n_2944), .A1 (inputB[13]), .A2 (inputA[14]));
NOR3_X1 i_3737 (.ZN (n_2943), .A1 (n_880), .A2 (n_2944), .A3 (n_529));
AOI22_X1 i_3736 (.ZN (n_2942), .A1 (inputB[12]), .A2 (inputA[14]), .B1 (inputB[13]), .B2 (inputA[13]));
NOR2_X1 i_3735 (.ZN (n_2941), .A1 (n_2943), .A2 (n_2942));
NAND2_X1 i_3734 (.ZN (n_2940), .A1 (inputB[14]), .A2 (inputA[12]));
INV_X1 i_3733 (.ZN (n_2939), .A (n_2940));
AOI21_X1 i_3732 (.ZN (n_2938), .A (n_2943), .B1 (n_2941), .B2 (n_2939));
OAI21_X1 i_3731 (.ZN (n_2937), .A (n_2946), .B1 (n_2945), .B2 (n_2938));
XNOR2_X1 i_3730 (.ZN (n_2936), .A (n_2960), .B (n_2937));
NAND2_X1 i_3729 (.ZN (n_2935), .A1 (inputB[2]), .A2 (inputA[25]));
XNOR2_X1 i_3728 (.ZN (n_2934), .A (n_2998), .B (n_2935));
NAND2_X1 i_3727 (.ZN (n_2933), .A1 (inputB[3]), .A2 (inputA[24]));
OAI22_X1 i_3726 (.ZN (n_2932), .A1 (n_2998), .A2 (n_2935), .B1 (n_2934), .B2 (n_2933));
NOR2_X1 i_3725 (.ZN (n_2931), .A1 (n_215), .A2 (n_63));
XOR2_X1 i_3724 (.Z (n_2930), .A (n_2932), .B (n_2931));
NAND2_X1 i_3723 (.ZN (n_2929), .A1 (inputB[0]), .A2 (inputA[28]));
XOR2_X1 i_3722 (.Z (n_2928), .A (n_2930), .B (n_2929));
XNOR2_X1 i_3721 (.ZN (n_2927), .A (n_2936), .B (n_2928));
NAND2_X1 i_3720 (.ZN (n_2926), .A1 (inputB[1]), .A2 (inputA[23]));
NAND2_X1 i_3719 (.ZN (n_2925), .A1 (inputB[2]), .A2 (inputA[22]));
XNOR2_X1 i_3718 (.ZN (n_2924), .A (n_2926), .B (n_2925));
NAND2_X1 i_3717 (.ZN (n_2923), .A1 (inputB[3]), .A2 (inputA[21]));
AOI22_X1 i_3716 (.ZN (n_2911), .A1 (n_2670), .A2 (n_2666), .B1 (n_2665), .B2 (n_2658));
AOI22_X1 i_3715 (.ZN (n_2910), .A1 (n_2646), .A2 (n_2649), .B1 (n_2645), .B2 (n_2653));
INV_X1 i_3714 (.ZN (n_2909), .A (n_2910));
XOR2_X1 i_3713 (.Z (n_2908), .A (n_2924), .B (n_2923));
XOR2_X1 i_3712 (.Z (n_2907), .A (n_2909), .B (n_2908));
NAND2_X1 i_3711 (.ZN (n_2904), .A1 (n_2911), .A2 (n_2907));
OAI21_X1 i_3710 (.ZN (n_2903), .A (n_2904), .B1 (n_2911), .B2 (n_2907));
NOR2_X1 i_3709 (.ZN (n_2902), .A1 (n_2691), .A2 (n_2926));
AOI22_X1 i_3708 (.ZN (n_2901), .A1 (inputB[0]), .A2 (inputA[23]), .B1 (inputB[1]), .B2 (inputA[22]));
NOR2_X1 i_3707 (.ZN (n_2900), .A1 (n_2902), .A2 (n_2901));
NOR2_X1 i_3705 (.ZN (n_2899), .A1 (n_1219), .A2 (n_482));
OAI21_X1 i_3703 (.ZN (n_2898), .A (n_2688), .B1 (n_2689), .B2 (n_2687));
INV_X1 i_3702 (.ZN (n_2896), .A (n_2898));
XOR2_X1 i_3701 (.Z (n_2895), .A (n_2900), .B (n_2899));
XOR2_X1 i_3700 (.Z (n_2894), .A (n_2896), .B (n_2895));
NAND2_X1 i_3699 (.ZN (n_2891), .A1 (inputB[4]), .A2 (inputA[20]));
NOR2_X1 i_3698 (.ZN (n_2890), .A1 (n_2669), .A2 (n_2891));
AOI22_X1 i_3696 (.ZN (n_2889), .A1 (inputB[3]), .A2 (inputA[20]), .B1 (inputB[4]), .B2 (inputA[19]));
NOR2_X1 i_3695 (.ZN (n_2888), .A1 (n_2890), .A2 (n_2889));
NOR2_X1 i_3694 (.ZN (n_2887), .A1 (n_668), .A2 (n_479));
XOR2_X1 i_3693 (.Z (n_2884), .A (n_2888), .B (n_2887));
OAI21_X1 i_3692 (.ZN (n_2883), .A (n_2783), .B1 (n_2784), .B2 (n_2788));
XOR2_X1 i_3691 (.Z (n_2882), .A (n_2775), .B (n_2774));
XOR2_X1 i_3690 (.Z (n_2880), .A (n_2883), .B (n_2882));
XNOR2_X1 i_3689 (.ZN (n_2879), .A (n_2767), .B (n_2766));
AOI22_X1 i_3688 (.ZN (n_2877), .A1 (n_2883), .A2 (n_2882), .B1 (n_2880), .B2 (n_2879));
INV_X1 i_3687 (.ZN (n_2876), .A (n_2877));
AOI22_X1 i_3686 (.ZN (n_2875), .A1 (n_2896), .A2 (n_2895), .B1 (n_2894), .B2 (n_2884));
NOR2_X1 i_3685 (.ZN (n_2874), .A1 (n_2876), .A2 (n_2875));
AOI21_X1 i_3684 (.ZN (n_2873), .A (n_2874), .B1 (n_2876), .B2 (n_2875));
AOI21_X1 i_3683 (.ZN (n_2851), .A (n_2874), .B1 (n_2903), .B2 (n_2873));
NAND2_X1 i_3682 (.ZN (n_2850), .A1 (inputB[14]), .A2 (inputA[10]));
NAND2_X1 i_3681 (.ZN (n_2849), .A1 (inputB[17]), .A2 (inputA[8]));
NAND2_X1 i_3680 (.ZN (n_2848), .A1 (inputB[18]), .A2 (inputA[6]));
XNOR2_X1 i_3679 (.ZN (n_2847), .A (n_2770), .B (n_2850));
NAND2_X1 i_3678 (.ZN (n_2846), .A1 (inputB[15]), .A2 (inputA[9]));
OAI22_X1 i_3677 (.ZN (n_2845), .A1 (n_2770), .A2 (n_2850), .B1 (n_2847), .B2 (n_2846));
NOR2_X1 i_3676 (.ZN (n_2844), .A1 (n_2753), .A2 (n_2849));
AOI22_X1 i_3675 (.ZN (n_2843), .A1 (inputB[16]), .A2 (inputA[8]), .B1 (inputB[17]), .B2 (inputA[7]));
OR2_X1 i_3674 (.ZN (n_2842), .A1 (n_2844), .A2 (n_2843));
NOR2_X1 i_3673 (.ZN (n_2841), .A1 (n_2848), .A2 (n_2842));
OR2_X1 i_3672 (.ZN (n_2840), .A1 (n_2844), .A2 (n_2841));
NAND2_X1 i_3671 (.ZN (n_2839), .A1 (n_2845), .A2 (n_2840));
OAI21_X1 i_3670 (.ZN (n_2838), .A (n_2839), .B1 (n_2845), .B2 (n_2840));
NAND2_X1 i_3669 (.ZN (n_2837), .A1 (inputB[20]), .A2 (inputA[4]));
XNOR2_X1 i_3668 (.ZN (n_2836), .A (n_2749), .B (n_2837));
NAND2_X1 i_3667 (.ZN (n_2835), .A1 (inputB[21]), .A2 (inputA[3]));
OAI22_X1 i_3666 (.ZN (n_2834), .A1 (n_2749), .A2 (n_2837), .B1 (n_2836), .B2 (n_2835));
XOR2_X1 i_3665 (.Z (n_2833), .A (n_2838), .B (n_2834));
INV_X1 i_3664 (.ZN (n_2831), .A (n_2833));
NAND2_X1 i_3663 (.ZN (n_2830), .A1 (inputB[23]), .A2 (inputA[2]));
XNOR2_X1 i_3662 (.ZN (n_2829), .A (n_2763), .B (n_2830));
NAND2_X1 i_3661 (.ZN (n_2828), .A1 (inputB[25]), .A2 (inputA[0]));
XOR2_X1 i_3660 (.Z (n_2826), .A (n_2829), .B (n_2828));
XNOR2_X1 i_3659 (.ZN (n_2825), .A (n_2833), .B (n_2826));
NAND2_X1 i_3658 (.ZN (n_2824), .A1 (inputB[9]), .A2 (inputA[16]));
AOI22_X1 i_3657 (.ZN (n_2823), .A1 (inputB[8]), .A2 (inputA[16]), .B1 (inputB[9]), .B2 (inputA[15]));
INV_X1 i_3656 (.ZN (n_2822), .A (n_2823));
OAI21_X1 i_3655 (.ZN (n_2821), .A (n_2822), .B1 (n_2774), .B2 (n_2824));
OAI22_X1 i_3654 (.ZN (n_2820), .A1 (n_2774), .A2 (n_2824), .B1 (n_2782), .B2 (n_2821));
INV_X1 i_3653 (.ZN (n_2819), .A (n_2820));
NAND2_X1 i_3652 (.ZN (n_2818), .A1 (inputB[5]), .A2 (inputA[19]));
XNOR2_X1 i_3651 (.ZN (n_2817), .A (n_2891), .B (n_2818));
NAND2_X1 i_3650 (.ZN (n_2816), .A1 (inputB[6]), .A2 (inputA[18]));
OAI22_X1 i_3649 (.ZN (n_2815), .A1 (n_2891), .A2 (n_2818), .B1 (n_2817), .B2 (n_2816));
XOR2_X1 i_3648 (.Z (n_2814), .A (n_2819), .B (n_2815));
OR2_X1 i_3647 (.ZN (n_2813), .A1 (n_1131), .A2 (n_530));
OR2_X1 i_3646 (.ZN (n_2812), .A1 (n_667), .A2 (n_880));
XNOR2_X1 i_3645 (.ZN (n_2811), .A (n_2787), .B (n_2813));
OAI22_X1 i_3644 (.ZN (n_2810), .A1 (n_2787), .A2 (n_2813), .B1 (n_2812), .B2 (n_2811));
INV_X1 i_3643 (.ZN (n_2809), .A (n_2810));
XOR2_X1 i_3642 (.Z (n_2808), .A (n_2814), .B (n_2809));
XNOR2_X1 i_3641 (.ZN (n_2807), .A (n_2825), .B (n_2808));
XOR2_X1 i_3640 (.Z (n_2806), .A (n_2851), .B (n_2807));
OAI21_X1 i_3639 (.ZN (n_2805), .A (n_2904), .B1 (n_2909), .B2 (n_2908));
INV_X1 i_3638 (.ZN (n_2804), .A (n_2805));
XOR2_X1 i_3637 (.Z (n_2803), .A (n_2817), .B (n_2816));
XOR2_X1 i_3636 (.Z (n_2802), .A (n_2782), .B (n_2821));
NOR2_X1 i_3635 (.ZN (n_2801), .A1 (n_2803), .A2 (n_2802));
AOI21_X1 i_3634 (.ZN (n_2800), .A (n_2801), .B1 (n_2803), .B2 (n_2802));
XNOR2_X1 i_3633 (.ZN (n_2799), .A (n_2812), .B (n_2811));
AOI21_X1 i_3632 (.ZN (n_2798), .A (n_2801), .B1 (n_2800), .B2 (n_2799));
AOI21_X1 i_3631 (.ZN (n_2797), .A (n_2841), .B1 (n_2848), .B2 (n_2842));
XOR2_X1 i_3630 (.Z (n_2796), .A (n_2847), .B (n_2846));
NOR2_X1 i_3629 (.ZN (n_2795), .A1 (n_2797), .A2 (n_2796));
AOI21_X1 i_3628 (.ZN (n_2794), .A (n_2795), .B1 (n_2797), .B2 (n_2796));
XNOR2_X1 i_3627 (.ZN (n_2793), .A (n_2836), .B (n_2835));
AOI21_X1 i_3626 (.ZN (n_2792), .A (n_2795), .B1 (n_2794), .B2 (n_2793));
XOR2_X1 i_3625 (.Z (n_2791), .A (n_2798), .B (n_2792));
XOR2_X1 i_3624 (.Z (n_2790), .A (n_2805), .B (n_2791));
XNOR2_X1 i_3623 (.ZN (n_2789), .A (n_2806), .B (n_2790));
INV_X1 i_3622 (.ZN (n_2788), .A (n_2664));
NAND2_X1 i_3621 (.ZN (n_2787), .A1 (inputB[11]), .A2 (inputA[13]));
NOR2_X1 i_3620 (.ZN (n_2786), .A1 (n_2659), .A2 (n_2787));
AOI22_X1 i_3619 (.ZN (n_2785), .A1 (inputB[10]), .A2 (inputA[13]), .B1 (inputB[11]), .B2 (inputA[12]));
NOR2_X1 i_3618 (.ZN (n_2784), .A1 (n_2786), .A2 (n_2785));
NAND2_X1 i_3617 (.ZN (n_2783), .A1 (n_2788), .A2 (n_2784));
NAND2_X1 i_3616 (.ZN (n_2782), .A1 (inputB[7]), .A2 (inputA[17]));
NOR2_X1 i_3615 (.ZN (n_2777), .A1 (n_2674), .A2 (n_2782));
AOI22_X1 i_3614 (.ZN (n_2776), .A1 (inputB[7]), .A2 (inputA[16]), .B1 (inputB[6]), .B2 (inputA[17]));
NOR2_X1 i_3613 (.ZN (n_2775), .A1 (n_2777), .A2 (n_2776));
NAND2_X1 i_3612 (.ZN (n_2774), .A1 (inputB[8]), .A2 (inputA[15]));
OAI21_X1 i_3611 (.ZN (n_2773), .A (n_2783), .B1 (n_2659), .B2 (n_2787));
OAI22_X1 i_3610 (.ZN (n_2772), .A1 (n_2674), .A2 (n_2782), .B1 (n_2776), .B2 (n_2774));
XOR2_X1 i_3609 (.Z (n_2771), .A (n_2773), .B (n_2772));
NAND2_X1 i_3608 (.ZN (n_2770), .A1 (inputB[13]), .A2 (inputA[11]));
AOI22_X1 i_3607 (.ZN (n_2769), .A1 (inputB[13]), .A2 (inputA[10]), .B1 (inputB[12]), .B2 (inputA[11]));
INV_X1 i_3606 (.ZN (n_2768), .A (n_2769));
OAI21_X1 i_3605 (.ZN (n_2767), .A (n_2768), .B1 (n_2621), .B2 (n_2770));
NAND2_X1 i_3604 (.ZN (n_2766), .A1 (inputB[14]), .A2 (inputA[9]));
OAI22_X1 i_3603 (.ZN (n_2765), .A1 (n_2621), .A2 (n_2770), .B1 (n_2767), .B2 (n_2766));
NAND2_X1 i_3602 (.ZN (n_2764), .A1 (inputB[23]), .A2 (inputA[0]));
NAND2_X1 i_3601 (.ZN (n_2763), .A1 (inputB[24]), .A2 (inputA[1]));
NOR2_X1 i_3599 (.ZN (n_2762), .A1 (n_2764), .A2 (n_2763));
AOI22_X1 i_3598 (.ZN (n_2761), .A1 (inputB[23]), .A2 (inputA[1]), .B1 (inputB[24]), .B2 (inputA[0]));
NOR2_X1 i_3597 (.ZN (n_2760), .A1 (n_2762), .A2 (n_2761));
NAND2_X1 i_3596 (.ZN (n_2759), .A1 (inputB[22]), .A2 (inputA[2]));
INV_X1 i_3595 (.ZN (n_2758), .A (n_2759));
AOI21_X1 i_3594 (.ZN (n_2757), .A (n_2762), .B1 (n_2760), .B2 (n_2758));
AOI22_X1 i_3593 (.ZN (n_2756), .A1 (n_2773), .A2 (n_2772), .B1 (n_2771), .B2 (n_2765));
NAND2_X1 i_3592 (.ZN (n_2755), .A1 (n_2757), .A2 (n_2756));
OR2_X1 i_3591 (.ZN (n_2754), .A1 (n_2757), .A2 (n_2756));
NAND2_X1 i_3590 (.ZN (n_2753), .A1 (inputB[16]), .A2 (inputA[7]));
NAND2_X1 i_3589 (.ZN (n_2752), .A1 (inputB[15]), .A2 (inputA[8]));
XNOR2_X1 i_3588 (.ZN (n_2751), .A (n_2753), .B (n_2752));
NAND2_X1 i_3587 (.ZN (n_2750), .A1 (inputB[17]), .A2 (inputA[6]));
NAND2_X1 i_3586 (.ZN (n_2749), .A1 (inputB[19]), .A2 (inputA[5]));
NOR2_X1 i_3585 (.ZN (n_2748), .A1 (n_2655), .A2 (n_2749));
AOI22_X1 i_3584 (.ZN (n_2747), .A1 (inputB[19]), .A2 (inputA[4]), .B1 (inputB[18]), .B2 (inputA[5]));
NOR2_X1 i_3583 (.ZN (n_2746), .A1 (n_2748), .A2 (n_2747));
NOR2_X1 i_3582 (.ZN (n_2745), .A1 (n_1724), .A2 (n_414));
AOI21_X1 i_3581 (.ZN (n_2744), .A (n_2748), .B1 (n_2746), .B2 (n_2745));
INV_X1 i_3580 (.ZN (n_2743), .A (n_2744));
OAI22_X1 i_3579 (.ZN (n_2742), .A1 (n_2753), .A2 (n_2752), .B1 (n_2751), .B2 (n_2750));
XOR2_X1 i_3578 (.Z (n_2741), .A (n_2743), .B (n_2742));
NAND2_X1 i_3577 (.ZN (n_2740), .A1 (inputB[21]), .A2 (inputA[1]));
NOR2_X1 i_3576 (.ZN (n_2739), .A1 (n_2759), .A2 (n_2740));
INV_X1 i_3575 (.ZN (n_2738), .A (n_2739));
AOI22_X1 i_3574 (.ZN (n_2718), .A1 (inputB[22]), .A2 (inputA[1]), .B1 (inputB[21]), .B2 (inputA[2]));
NOR2_X1 i_3573 (.ZN (n_2717), .A1 (n_2739), .A2 (n_2718));
AOI21_X1 i_3572 (.ZN (n_2716), .A (n_2718), .B1 (n_2764), .B2 (n_2738));
INV_X1 i_3571 (.ZN (n_2715), .A (n_2716));
AOI22_X1 i_3570 (.ZN (n_2714), .A1 (n_2743), .A2 (n_2742), .B1 (n_2741), .B2 (n_2716));
NAND2_X1 i_3569 (.ZN (n_2713), .A1 (n_2754), .A2 (n_2714));
NAND2_X1 i_3568 (.ZN (n_2712), .A1 (n_2755), .A2 (n_2713));
NAND2_X1 i_3567 (.ZN (n_2711), .A1 (inputB[25]), .A2 (inputA[1]));
NAND2_X1 i_3566 (.ZN (n_2710), .A1 (inputB[26]), .A2 (inputA[0]));
XOR2_X1 i_3565 (.Z (n_2709), .A (n_2711), .B (n_2710));
INV_X1 i_3564 (.ZN (n_2708), .A (n_2709));
NAND2_X1 i_3563 (.ZN (n_2707), .A1 (inputB[24]), .A2 (inputA[2]));
XOR2_X1 i_3562 (.Z (n_2706), .A (n_2709), .B (n_2707));
NAND2_X1 i_3561 (.ZN (n_2705), .A1 (inputB[21]), .A2 (inputA[5]));
NAND2_X1 i_3560 (.ZN (n_2704), .A1 (inputB[22]), .A2 (inputA[4]));
XOR2_X1 i_3559 (.Z (n_2703), .A (n_2705), .B (n_2704));
INV_X1 i_3558 (.ZN (n_2702), .A (n_2703));
NAND2_X1 i_3557 (.ZN (n_2701), .A1 (inputB[23]), .A2 (inputA[3]));
XOR2_X1 i_3556 (.Z (n_2700), .A (n_2703), .B (n_2701));
XNOR2_X1 i_3555 (.ZN (n_2698), .A (n_2706), .B (n_2700));
XOR2_X1 i_3554 (.Z (n_2697), .A (n_2712), .B (n_2698));
OAI21_X1 i_3553 (.ZN (n_2696), .A (n_2542), .B1 (n_2532), .B2 (n_2534));
INV_X1 i_3552 (.ZN (n_2695), .A (n_2696));
AOI22_X1 i_3551 (.ZN (n_2694), .A1 (n_2544), .A2 (n_2546), .B1 (n_2547), .B2 (n_2548));
NOR2_X1 i_3550 (.ZN (n_2693), .A1 (n_2695), .A2 (n_2694));
AOI21_X1 i_3549 (.ZN (n_2692), .A (n_2693), .B1 (n_2695), .B2 (n_2694));
NAND2_X1 i_3548 (.ZN (n_2691), .A1 (inputB[0]), .A2 (inputA[22]));
AOI21_X1 i_3547 (.ZN (n_2690), .A (n_2600), .B1 (n_2598), .B2 (n_2597));
NOR2_X1 i_3546 (.ZN (n_2689), .A1 (n_2691), .A2 (n_2690));
NAND2_X1 i_3545 (.ZN (n_2688), .A1 (n_2691), .A2 (n_2690));
NOR2_X1 i_3544 (.ZN (n_2687), .A1 (n_63), .A2 (n_482));
AOI21_X1 i_3543 (.ZN (n_2686), .A (n_2689), .B1 (n_2691), .B2 (n_2690));
XOR2_X1 i_3542 (.Z (n_2685), .A (n_2687), .B (n_2686));
XOR2_X1 i_3541 (.Z (n_2684), .A (n_2660), .B (n_2659));
XOR2_X1 i_3540 (.Z (n_2683), .A (n_2668), .B (n_2667));
XOR2_X1 i_3539 (.Z (n_2681), .A (n_2684), .B (n_2683));
XNOR2_X1 i_3538 (.ZN (n_2680), .A (n_2672), .B (n_2671));
NAND2_X1 i_3537 (.ZN (n_2679), .A1 (n_2681), .A2 (n_2680));
OAI21_X1 i_3536 (.ZN (n_2678), .A (n_2679), .B1 (n_2684), .B2 (n_2683));
AOI21_X1 i_3535 (.ZN (n_2677), .A (n_2693), .B1 (n_2692), .B2 (n_2685));
NAND2_X1 i_3534 (.ZN (n_2676), .A1 (n_2678), .A2 (n_2677));
OAI21_X1 i_3533 (.ZN (n_2675), .A (n_2676), .B1 (n_2678), .B2 (n_2677));
NAND2_X1 i_3532 (.ZN (n_2674), .A1 (inputB[6]), .A2 (inputA[16]));
NAND2_X1 i_3531 (.ZN (n_2673), .A1 (inputB[5]), .A2 (inputA[17]));
XNOR2_X1 i_3530 (.ZN (n_2672), .A (n_2674), .B (n_2673));
NAND2_X1 i_3529 (.ZN (n_2671), .A1 (inputB[7]), .A2 (inputA[15]));
OAI22_X1 i_3528 (.ZN (n_2670), .A1 (n_2674), .A2 (n_2673), .B1 (n_2672), .B2 (n_2671));
NAND2_X1 i_3527 (.ZN (n_2669), .A1 (inputB[3]), .A2 (inputA[19]));
XNOR2_X1 i_3526 (.ZN (n_2668), .A (n_2601), .B (n_2669));
NAND2_X1 i_3525 (.ZN (n_2667), .A1 (inputB[4]), .A2 (inputA[18]));
OAI22_X1 i_3524 (.ZN (n_2666), .A1 (n_2601), .A2 (n_2669), .B1 (n_2668), .B2 (n_2667));
XOR2_X1 i_3523 (.Z (n_2665), .A (n_2670), .B (n_2666));
NAND2_X1 i_3522 (.ZN (n_2664), .A1 (inputB[9]), .A2 (inputA[14]));
AOI22_X1 i_3521 (.ZN (n_2662), .A1 (inputB[9]), .A2 (inputA[13]), .B1 (inputB[8]), .B2 (inputA[14]));
INV_X1 i_3520 (.ZN (n_2661), .A (n_2662));
OAI21_X1 i_3519 (.ZN (n_2660), .A (n_2661), .B1 (n_1964), .B2 (n_2664));
NAND2_X1 i_3518 (.ZN (n_2659), .A1 (inputB[10]), .A2 (inputA[12]));
OAI22_X1 i_3517 (.ZN (n_2658), .A1 (n_1964), .A2 (n_2664), .B1 (n_2660), .B2 (n_2659));
XOR2_X1 i_3516 (.Z (n_2657), .A (n_2665), .B (n_2658));
NAND2_X1 i_3515 (.ZN (n_2656), .A1 (inputB[17]), .A2 (inputA[5]));
NAND2_X1 i_3514 (.ZN (n_2655), .A1 (inputB[18]), .A2 (inputA[4]));
XNOR2_X1 i_3513 (.ZN (n_2654), .A (n_2656), .B (n_2655));
OAI33_X1 i_3512 (.ZN (n_2653), .A1 (n_1724), .A2 (n_314), .A3 (n_2654), .B1 (n_859)
    , .B2 (n_881), .B3 (n_2655));
NAND2_X1 i_3511 (.ZN (n_2652), .A1 (inputB[15]), .A2 (inputA[7]));
XNOR2_X1 i_3510 (.ZN (n_2651), .A (n_2634), .B (n_2652));
NAND2_X1 i_3509 (.ZN (n_2650), .A1 (inputB[16]), .A2 (inputA[6]));
OAI22_X1 i_3508 (.ZN (n_2649), .A1 (n_2634), .A2 (n_2652), .B1 (n_2651), .B2 (n_2650));
NAND2_X1 i_3507 (.ZN (n_2648), .A1 (inputB[11]), .A2 (inputA[11]));
XNOR2_X1 i_3506 (.ZN (n_2647), .A (n_2621), .B (n_2648));
OAI33_X1 i_3505 (.ZN (n_2646), .A1 (n_1894), .A2 (n_671), .A3 (n_2647), .B1 (n_2621)
    , .B2 (n_670), .B3 (n_1136));
XOR2_X1 i_3504 (.Z (n_2645), .A (n_2649), .B (n_2646));
XOR2_X1 i_3503 (.Z (n_2636), .A (n_2653), .B (n_2645));
XOR2_X1 i_3502 (.Z (n_2635), .A (n_2657), .B (n_2636));
NAND2_X1 i_3501 (.ZN (n_2634), .A1 (inputB[14]), .A2 (inputA[8]));
NOR2_X1 i_3500 (.ZN (n_2633), .A1 (n_2530), .A2 (n_2634));
AOI22_X1 i_3499 (.ZN (n_2632), .A1 (inputB[13]), .A2 (inputA[8]), .B1 (inputB[14]), .B2 (inputA[7]));
NOR2_X1 i_3498 (.ZN (n_2630), .A1 (n_2633), .A2 (n_2632));
NOR2_X1 i_3497 (.ZN (n_2629), .A1 (n_1349), .A2 (n_587));
NAND2_X1 i_3496 (.ZN (n_2628), .A1 (inputB[7]), .A2 (inputA[14]));
XOR2_X1 i_3495 (.Z (n_2627), .A (n_1964), .B (n_2628));
AND2_X1 i_3494 (.ZN (n_2626), .A1 (inputB[9]), .A2 (inputA[12]));
NAND2_X1 i_3493 (.ZN (n_2625), .A1 (n_2627), .A2 (n_2626));
OAI21_X1 i_3492 (.ZN (n_2624), .A (n_2625), .B1 (n_2627), .B2 (n_2626));
XNOR2_X1 i_3491 (.ZN (n_2623), .A (n_2630), .B (n_2629));
XOR2_X1 i_3490 (.Z (n_2622), .A (n_2624), .B (n_2623));
NAND2_X1 i_3489 (.ZN (n_2621), .A1 (inputB[12]), .A2 (inputA[10]));
NOR2_X1 i_3488 (.ZN (n_2620), .A1 (n_1934), .A2 (n_2621));
AOI22_X1 i_3487 (.ZN (n_2619), .A1 (inputB[12]), .A2 (inputA[9]), .B1 (inputB[11]), .B2 (inputA[10]));
OR2_X1 i_3485 (.ZN (n_2618), .A1 (n_2620), .A2 (n_2619));
NOR2_X1 i_3484 (.ZN (n_2617), .A1 (n_1938), .A2 (n_2618));
AOI21_X1 i_3483 (.ZN (n_2616), .A (n_2617), .B1 (n_1938), .B2 (n_2618));
INV_X1 i_3482 (.ZN (n_2615), .A (n_2616));
AOI22_X1 i_3481 (.ZN (n_2613), .A1 (n_2624), .A2 (n_2623), .B1 (n_2622), .B2 (n_2615));
OAI21_X1 i_3480 (.ZN (n_2612), .A (n_2625), .B1 (n_1964), .B2 (n_2628));
OR2_X1 i_3479 (.ZN (n_2611), .A1 (n_668), .A2 (n_865));
NAND2_X1 i_3478 (.ZN (n_2610), .A1 (n_1948), .A2 (n_2611));
NOR2_X1 i_3477 (.ZN (n_2609), .A1 (n_1948), .A2 (n_2611));
NOR2_X1 i_3476 (.ZN (n_2608), .A1 (n_878), .A2 (n_478));
OAI21_X1 i_3475 (.ZN (n_2607), .A (n_2610), .B1 (n_2609), .B2 (n_2608));
XNOR2_X1 i_3474 (.ZN (n_2606), .A (n_2612), .B (n_2607));
NOR2_X1 i_3473 (.ZN (n_2605), .A1 (n_2620), .A2 (n_2617));
INV_X1 i_3472 (.ZN (n_2604), .A (n_2605));
XOR2_X1 i_3471 (.Z (n_2603), .A (n_2606), .B (n_2605));
XNOR2_X1 i_3470 (.ZN (n_2602), .A (n_2613), .B (n_2603));
NAND2_X1 i_3469 (.ZN (n_2601), .A1 (inputB[2]), .A2 (inputA[20]));
NOR2_X1 i_3468 (.ZN (n_2600), .A1 (n_2013), .A2 (n_2601));
AOI22_X1 i_3467 (.ZN (n_2599), .A1 (inputB[1]), .A2 (inputA[20]), .B1 (inputB[2]), .B2 (inputA[19]));
NOR2_X1 i_3466 (.ZN (n_2598), .A1 (n_2600), .A2 (n_2599));
NOR2_X1 i_3465 (.ZN (n_2597), .A1 (n_685), .A2 (n_479));
NAND2_X1 i_3464 (.ZN (n_2590), .A1 (n_1923), .A2 (n_1928));
OAI21_X1 i_3463 (.ZN (n_2589), .A (n_2590), .B1 (n_1914), .B2 (n_1922));
XOR2_X1 i_3462 (.Z (n_2588), .A (n_2598), .B (n_2597));
XOR2_X1 i_3461 (.Z (n_2587), .A (n_2589), .B (n_2588));
OAI21_X1 i_3460 (.ZN (n_2586), .A (n_2610), .B1 (n_1948), .B2 (n_2611));
XNOR2_X1 i_3459 (.ZN (n_2585), .A (n_2608), .B (n_2586));
AOI22_X1 i_3458 (.ZN (n_2584), .A1 (n_2589), .A2 (n_2588), .B1 (n_2587), .B2 (n_2585));
XNOR2_X1 i_3457 (.ZN (n_2583), .A (n_2602), .B (n_2584));
AOI22_X1 i_3456 (.ZN (n_2582), .A1 (n_2581), .A2 (n_2578), .B1 (n_2579), .B2 (n_2580));
XOR2_X1 i_3455 (.Z (n_2581), .A (n_2579), .B (n_2580));
AOI22_X1 i_3454 (.ZN (n_2580), .A1 (n_2003), .A2 (n_1995), .B1 (n_1994), .B2 (n_1966));
XNOR2_X1 i_3453 (.ZN (n_2579), .A (n_2550), .B (n_2565));
XOR2_X1 i_3452 (.Z (n_2578), .A (n_2566), .B (n_2577));
XOR2_X1 i_3451 (.Z (n_2577), .A (n_2574), .B (n_2576));
AOI22_X1 i_3450 (.ZN (n_2576), .A1 (n_1940), .A2 (n_1960), .B1 (n_1939), .B2 (n_1933));
AOI22_X1 i_3449 (.ZN (n_2574), .A1 (n_2573), .A2 (n_1974), .B1 (n_1972), .B2 (n_1967));
INV_X1 i_3448 (.ZN (n_2573), .A (n_1973));
AOI22_X1 i_3447 (.ZN (n_2566), .A1 (n_1895), .A2 (n_1904), .B1 (n_1905), .B2 (n_1929));
OAI21_X1 i_3446 (.ZN (n_2565), .A (n_2557), .B1 (n_2558), .B2 (n_2564));
XOR2_X1 i_3445 (.Z (n_2564), .A (n_2562), .B (n_2563));
NAND2_X1 i_3444 (.ZN (n_2563), .A1 (inputA[0]), .A2 (inputB[20]));
NAND2_X1 i_3443 (.ZN (n_2562), .A1 (n_2560), .A2 (n_2561));
OAI22_X1 i_3442 (.ZN (n_2561), .A1 (n_314), .A2 (n_1547), .B1 (n_67), .B2 (n_400));
NAND3_X1 i_3441 (.ZN (n_2560), .A1 (n_2559), .A2 (inputA[1]), .A3 (inputB[18]));
NOR2_X1 i_3440 (.ZN (n_2559), .A1 (n_314), .A2 (n_67));
NOR2_X1 i_3439 (.ZN (n_2558), .A1 (n_2554), .A2 (n_2556));
NAND2_X1 i_3438 (.ZN (n_2557), .A1 (n_2554), .A2 (n_2556));
XNOR2_X1 i_3437 (.ZN (n_2556), .A (n_2555), .B (n_2552));
XNOR2_X1 i_3436 (.ZN (n_2555), .A (n_2551), .B (n_1723));
XNOR2_X1 i_3435 (.ZN (n_2554), .A (n_2539), .B (n_2553));
NAND2_X1 i_3434 (.ZN (n_2553), .A1 (inputA[6]), .A2 (inputB[14]));
NAND2_X1 i_3433 (.ZN (n_2552), .A1 (inputA[3]), .A2 (inputB[17]));
NAND2_X1 i_3432 (.ZN (n_2551), .A1 (inputA[4]), .A2 (inputB[16]));
XOR2_X1 i_3431 (.Z (n_2550), .A (n_2543), .B (n_2549));
XNOR2_X1 i_3430 (.ZN (n_2549), .A (n_2547), .B (n_2548));
NOR2_X1 i_3429 (.ZN (n_2548), .A1 (n_62), .A2 (n_482));
XNOR2_X1 i_3428 (.ZN (n_2547), .A (n_2544), .B (n_2545));
INV_X1 i_3427 (.ZN (n_2546), .A (n_2545));
AOI21_X1 i_3426 (.ZN (n_2545), .A (n_1947), .B1 (n_1945), .B2 (n_1944));
OAI22_X1 i_3425 (.ZN (n_2544), .A1 (n_1969), .A2 (n_1968), .B1 (n_2013), .B2 (n_1971));
OAI21_X1 i_3424 (.ZN (n_2543), .A (n_2542), .B1 (n_2540), .B2 (n_2541));
NAND2_X1 i_3423 (.ZN (n_2542), .A1 (n_2540), .A2 (n_2541));
XOR2_X1 i_3422 (.Z (n_2541), .A (n_2532), .B (n_2534));
OAI33_X1 i_3421 (.ZN (n_2540), .A1 (n_2539), .A2 (n_1349), .A3 (n_586), .B1 (n_1898)
    , .B2 (n_1551), .B3 (n_671));
XNOR2_X1 i_3420 (.ZN (n_2539), .A (n_2530), .B (n_2535));
NAND2_X1 i_3419 (.ZN (n_2535), .A1 (inputA[8]), .A2 (inputB[12]));
AOI21_X1 i_3418 (.ZN (n_2534), .A (n_1937), .B1 (n_2533), .B2 (n_1935));
INV_X1 i_3417 (.ZN (n_2533), .A (n_1934));
AOI21_X1 i_3416 (.ZN (n_2532), .A (n_1963), .B1 (n_2531), .B2 (n_1961));
INV_X1 i_3415 (.ZN (n_2531), .A (n_1908));
NAND2_X1 i_3414 (.ZN (n_2530), .A1 (inputA[7]), .A2 (inputB[13]));
INV_X1 i_3413 (.ZN (n_2529), .A (n_2194));
XNOR2_X1 i_3412 (.ZN (n_2528), .A (n_2141), .B (n_2109));
XOR2_X1 i_3411 (.Z (n_2527), .A (n_2042), .B (n_2041));
NAND2_X1 i_3410 (.ZN (n_2526), .A1 (n_2528), .A2 (n_2527));
NOR2_X1 i_3409 (.ZN (n_2525), .A1 (n_2528), .A2 (n_2527));
AOI21_X1 i_3408 (.ZN (n_2524), .A (n_2525), .B1 (n_2528), .B2 (n_2527));
NOR3_X1 i_3407 (.ZN (n_2523), .A1 (n_2118), .A2 (n_529), .A3 (n_62));
INV_X1 i_3406 (.ZN (n_2522), .A (n_2523));
OAI22_X1 i_3405 (.ZN (n_2521), .A1 (n_529), .A2 (n_63), .B1 (n_62), .B2 (n_530));
NAND2_X1 i_3404 (.ZN (n_2520), .A1 (n_2522), .A2 (n_2521));
NAND2_X1 i_3403 (.ZN (n_2519), .A1 (inputB[2]), .A2 (inputA[12]));
NOR2_X1 i_3402 (.ZN (n_2518), .A1 (n_2520), .A2 (n_2519));
AOI21_X1 i_3401 (.ZN (n_2517), .A (n_2518), .B1 (n_2520), .B2 (n_2519));
NOR2_X1 i_3400 (.ZN (n_2513), .A1 (n_2134), .A2 (n_1844));
AOI21_X1 i_3399 (.ZN (n_2512), .A (n_2513), .B1 (n_2134), .B2 (n_1844));
INV_X1 i_3398 (.ZN (n_2511), .A (n_2512));
NAND2_X1 i_3397 (.ZN (n_2510), .A1 (inputB[5]), .A2 (inputA[9]));
NOR2_X1 i_3396 (.ZN (n_2509), .A1 (n_2511), .A2 (n_2510));
AOI21_X1 i_3395 (.ZN (n_2508), .A (n_2509), .B1 (n_2511), .B2 (n_2510));
NOR2_X1 i_3394 (.ZN (n_2507), .A1 (n_2517), .A2 (n_2508));
AOI21_X1 i_3393 (.ZN (n_2506), .A (n_2507), .B1 (n_2517), .B2 (n_2508));
NAND2_X1 i_3392 (.ZN (n_2505), .A1 (inputB[6]), .A2 (inputA[8]));
XNOR2_X1 i_3391 (.ZN (n_2504), .A (n_1843), .B (n_2505));
NAND2_X1 i_3390 (.ZN (n_2503), .A1 (inputB[8]), .A2 (inputA[6]));
XNOR2_X1 i_3389 (.ZN (n_2502), .A (n_2504), .B (n_2503));
XOR2_X1 i_3388 (.Z (n_2501), .A (n_2126), .B (n_2120));
NAND2_X1 i_3387 (.ZN (n_2500), .A1 (inputB[12]), .A2 (inputA[1]));
NOR2_X1 i_3386 (.ZN (n_2499), .A1 (n_16), .A2 (n_2500));
AOI22_X1 i_3385 (.ZN (n_2498), .A1 (inputB[13]), .A2 (inputA[1]), .B1 (inputB[12]), .B2 (inputA[2]));
NOR2_X1 i_3384 (.ZN (n_2497), .A1 (n_2499), .A2 (n_2498));
NOR2_X1 i_3383 (.ZN (n_2496), .A1 (n_66), .A2 (n_586));
XOR2_X1 i_3382 (.Z (n_2495), .A (n_2497), .B (n_2496));
AOI22_X1 i_3380 (.ZN (n_2494), .A1 (inputB[9]), .A2 (inputA[5]), .B1 (inputB[10]), .B2 (inputA[4]));
INV_X1 i_3379 (.ZN (n_2493), .A (n_2494));
OAI21_X1 i_3378 (.ZN (n_2492), .A (n_2493), .B1 (n_2125), .B2 (n_1828));
XOR2_X1 i_3377 (.Z (n_2491), .A (n_1833), .B (n_2492));
XOR2_X1 i_3376 (.Z (n_2489), .A (n_2495), .B (n_2491));
AOI21_X1 i_3375 (.ZN (n_2488), .A (n_2507), .B1 (n_2506), .B2 (n_2502));
INV_X1 i_3374 (.ZN (n_2487), .A (n_2488));
AOI22_X1 i_3373 (.ZN (n_2486), .A1 (n_2495), .A2 (n_2491), .B1 (n_2501), .B2 (n_2489));
NOR2_X1 i_3372 (.ZN (n_2485), .A1 (n_2487), .A2 (n_2486));
AOI21_X1 i_3371 (.ZN (n_2484), .A (n_2485), .B1 (n_2487), .B2 (n_2486));
XNOR2_X1 i_3370 (.ZN (n_2483), .A (n_2165), .B (n_2161));
AOI21_X1 i_3369 (.ZN (n_2482), .A (n_2485), .B1 (n_2484), .B2 (n_2483));
AOI21_X1 i_3368 (.ZN (n_2481), .A (n_2525), .B1 (n_2526), .B2 (n_2482));
XNOR2_X1 i_3367 (.ZN (n_2480), .A (n_2105), .B (n_2093));
NAND2_X1 i_3366 (.ZN (n_2479), .A1 (n_2481), .A2 (n_2480));
OAI21_X1 i_3365 (.ZN (n_2478), .A (n_2479), .B1 (n_2481), .B2 (n_2480));
XOR2_X1 i_3364 (.Z (n_2477), .A (n_1825), .B (n_1807));
XOR2_X1 i_3363 (.Z (n_2476), .A (n_2080), .B (n_2079));
XOR2_X1 i_3362 (.Z (n_2475), .A (n_2477), .B (n_2476));
OAI22_X1 i_3361 (.ZN (n_2473), .A1 (n_2125), .A2 (n_1828), .B1 (n_1833), .B2 (n_2492));
INV_X1 i_3360 (.ZN (n_2472), .A (n_2473));
OAI33_X1 i_3359 (.ZN (n_2471), .A1 (n_1349), .A2 (n_669), .A3 (n_2504), .B1 (n_1843)
    , .B2 (n_878), .B3 (n_1551));
INV_X1 i_3358 (.ZN (n_2470), .A (n_2471));
AOI21_X1 i_3357 (.ZN (n_2469), .A (n_2499), .B1 (n_2497), .B2 (n_2496));
OAI22_X1 i_3356 (.ZN (n_2468), .A1 (n_2472), .A2 (n_2470), .B1 (n_2473), .B2 (n_2471));
OAI22_X1 i_3355 (.ZN (n_2467), .A1 (n_2472), .A2 (n_2470), .B1 (n_2469), .B2 (n_2468));
OAI21_X1 i_3354 (.ZN (n_2466), .A (n_2164), .B1 (n_2163), .B2 (n_2162));
NOR2_X1 i_3353 (.ZN (n_2465), .A1 (n_2513), .A2 (n_2509));
NOR2_X1 i_3352 (.ZN (n_2464), .A1 (n_2523), .A2 (n_2518));
XNOR2_X1 i_3351 (.ZN (n_2463), .A (n_2104), .B (n_2465));
OAI22_X1 i_3350 (.ZN (n_2462), .A1 (n_2104), .A2 (n_2465), .B1 (n_2464), .B2 (n_2463));
XNOR2_X1 i_3349 (.ZN (n_2461), .A (n_2467), .B (n_2466));
OAI22_X1 i_3348 (.ZN (n_2460), .A1 (n_2467), .A2 (n_2466), .B1 (n_2462), .B2 (n_2461));
INV_X1 i_3347 (.ZN (n_2459), .A (n_2460));
XOR2_X1 i_3346 (.Z (n_2458), .A (n_2475), .B (n_2460));
XOR2_X1 i_3345 (.Z (n_2457), .A (n_2047), .B (n_2040));
XOR2_X1 i_3344 (.Z (n_2456), .A (n_2458), .B (n_2457));
XOR2_X1 i_3343 (.Z (n_2455), .A (n_2462), .B (n_2461));
XOR2_X1 i_3342 (.Z (n_2454), .A (n_2052), .B (n_2051));
XOR2_X1 i_3341 (.Z (n_2453), .A (n_2455), .B (n_2454));
NAND2_X1 i_3340 (.ZN (n_2452), .A1 (inputB[8]), .A2 (inputA[4]));
XNOR2_X1 i_3339 (.ZN (n_2451), .A (n_2202), .B (n_2452));
NAND2_X1 i_3338 (.ZN (n_2441), .A1 (inputB[9]), .A2 (inputA[3]));
NOR2_X1 i_3337 (.ZN (n_2440), .A1 (n_2185), .A2 (n_2136));
NOR2_X1 i_3336 (.ZN (n_2439), .A1 (n_15), .A2 (n_2440));
OAI22_X1 i_3335 (.ZN (n_2438), .A1 (n_2185), .A2 (n_2136), .B1 (n_15), .B2 (n_2140));
OAI22_X1 i_3334 (.ZN (n_2437), .A1 (n_2202), .A2 (n_2452), .B1 (n_2451), .B2 (n_2441));
XOR2_X1 i_3333 (.Z (n_2436), .A (n_2438), .B (n_2437));
NOR2_X1 i_3332 (.ZN (n_2435), .A1 (n_2189), .A2 (n_2500));
NOR2_X1 i_3331 (.ZN (n_2434), .A1 (n_14), .A2 (n_2435));
NAND2_X1 i_3330 (.ZN (n_2433), .A1 (n_2529), .A2 (n_2434));
OAI21_X1 i_3329 (.ZN (n_2432), .A (n_2433), .B1 (n_2189), .B2 (n_2500));
NAND2_X1 i_3328 (.ZN (n_2431), .A1 (inputB[11]), .A2 (inputA[2]));
XNOR2_X1 i_3327 (.ZN (n_2430), .A (n_2500), .B (n_2431));
NAND2_X1 i_3326 (.ZN (n_2429), .A1 (inputB[13]), .A2 (inputA[0]));
AOI22_X1 i_3325 (.ZN (n_2428), .A1 (n_2438), .A2 (n_2437), .B1 (n_2436), .B2 (n_2432));
INV_X1 i_3324 (.ZN (n_2427), .A (n_2428));
OAI22_X1 i_3323 (.ZN (n_2426), .A1 (n_2500), .A2 (n_2431), .B1 (n_2430), .B2 (n_2429));
NOR2_X1 i_3322 (.ZN (n_2425), .A1 (n_2427), .A2 (n_2426));
AOI21_X1 i_3321 (.ZN (n_2424), .A (n_2425), .B1 (n_2427), .B2 (n_2426));
AND3_X1 i_3320 (.ZN (n_2423), .A1 (inputB[1]), .A2 (n_2173), .A3 (inputA[13]));
XNOR2_X1 i_3319 (.ZN (n_2422), .A (n_2180), .B (n_2135));
OAI33_X1 i_3318 (.ZN (n_2421), .A1 (n_685), .A2 (n_1894), .A3 (n_2422), .B1 (n_63)
    , .B2 (n_2135), .B3 (n_1136));
AOI22_X1 i_3317 (.ZN (n_2420), .A1 (inputB[0]), .A2 (inputA[13]), .B1 (inputB[1]), .B2 (inputA[12]));
INV_X1 i_3316 (.ZN (n_2419), .A (n_2420));
AOI21_X1 i_3315 (.ZN (n_2418), .A (n_2423), .B1 (n_2421), .B2 (n_2419));
XOR2_X1 i_3314 (.Z (n_2417), .A (n_2469), .B (n_2468));
AOI21_X1 i_3313 (.ZN (n_2416), .A (n_2425), .B1 (n_2424), .B2 (n_2418));
XOR2_X1 i_3312 (.Z (n_2415), .A (n_2417), .B (n_2416));
XOR2_X1 i_3311 (.Z (n_2414), .A (n_2464), .B (n_2463));
AOI22_X1 i_3310 (.ZN (n_2413), .A1 (n_2417), .A2 (n_2416), .B1 (n_2415), .B2 (n_2414));
AOI22_X1 i_3309 (.ZN (n_2412), .A1 (n_2455), .A2 (n_2454), .B1 (n_2453), .B2 (n_2413));
XNOR2_X1 i_3308 (.ZN (n_2411), .A (n_2456), .B (n_2412));
OAI21_X1 i_3307 (.ZN (n_2410), .A (n_2479), .B1 (n_2478), .B2 (n_2411));
INV_X1 i_3306 (.ZN (n_2409), .A (n_10));
NOR2_X1 i_3305 (.ZN (n_2408), .A1 (n_62), .A2 (n_1349));
INV_X1 i_3304 (.ZN (n_2407), .A (n_2408));
XNOR2_X1 i_3303 (.ZN (n_2406), .A (n_2274), .B (n_13));
OAI33_X1 i_3302 (.ZN (n_2405), .A1 (n_1219), .A2 (n_1724), .A3 (n_2406), .B1 (n_62)
    , .B2 (n_2274), .B3 (n_859));
INV_X1 i_3301 (.ZN (n_2404), .A (n_2405));
XNOR2_X1 i_3300 (.ZN (n_2403), .A (n_9), .B (n_12));
NAND2_X1 i_3299 (.ZN (n_2402), .A1 (inputA[0]), .A2 (inputB[5]));
OAI22_X1 i_3298 (.ZN (n_2401), .A1 (n_9), .A2 (n_12), .B1 (n_2403), .B2 (n_2402));
INV_X1 i_3297 (.ZN (n_2400), .A (n_2401));
OAI22_X1 i_3296 (.ZN (n_2399), .A1 (n_2407), .A2 (n_2404), .B1 (n_2408), .B2 (n_2405));
OAI22_X1 i_3295 (.ZN (n_2398), .A1 (n_2407), .A2 (n_2404), .B1 (n_2400), .B2 (n_2399));
AOI22_X1 i_3294 (.ZN (n_2397), .A1 (inputA[1]), .A2 (inputB[5]), .B1 (inputA[2]), .B2 (inputB[4]));
INV_X1 i_3293 (.ZN (n_2396), .A (n_2397));
OAI21_X1 i_3292 (.ZN (n_2395), .A (n_2396), .B1 (n_12), .B2 (n_2279));
OAI22_X1 i_3291 (.ZN (n_2394), .A1 (n_12), .A2 (n_2279), .B1 (n_2283), .B2 (n_2395));
NAND2_X1 i_3290 (.ZN (n_2393), .A1 (n_2398), .A2 (n_2394));
OAI21_X1 i_3289 (.ZN (n_2392), .A (n_2393), .B1 (n_2398), .B2 (n_2394));
XOR2_X1 i_3288 (.Z (n_2385), .A (n_2269), .B (n_2266));
OAI21_X1 i_3287 (.ZN (n_2384), .A (n_2393), .B1 (n_2392), .B2 (n_2385));
XNOR2_X1 i_3286 (.ZN (n_2383), .A (n_2275), .B (n_2265));
NAND2_X1 i_3285 (.ZN (n_2382), .A1 (n_2384), .A2 (n_2383));
OAI21_X1 i_3284 (.ZN (n_2381), .A (n_2382), .B1 (n_2384), .B2 (n_2383));
XOR2_X1 i_3283 (.Z (n_2380), .A (n_2392), .B (n_2385));
XNOR2_X1 i_3282 (.ZN (n_2379), .A (n_2400), .B (n_2399));
XOR2_X1 i_3281 (.Z (n_2378), .A (n_2283), .B (n_2395));
XOR2_X1 i_3280 (.Z (n_2377), .A (n_2271), .B (n_2270));
NOR2_X1 i_3279 (.ZN (n_2376), .A1 (n_2378), .A2 (n_2377));
AOI21_X1 i_3278 (.ZN (n_2375), .A (n_2376), .B1 (n_2378), .B2 (n_2377));
AOI21_X1 i_3277 (.ZN (n_2374), .A (n_2376), .B1 (n_2379), .B2 (n_2375));
NAND2_X1 i_3276 (.ZN (n_2373), .A1 (n_2380), .A2 (n_2374));
OAI21_X1 i_3275 (.ZN (n_2372), .A (n_2382), .B1 (n_2381), .B2 (n_2373));
OAI33_X1 i_3274 (.ZN (n_2371), .A1 (n_76), .A2 (n_66), .A3 (n_685), .B1 (n_61), .B2 (n_63), .B3 (n_67));
AOI22_X1 i_3273 (.ZN (n_2370), .A1 (inputA[3]), .A2 (inputB[1]), .B1 (inputA[4]), .B2 (inputB[0]));
AOI21_X1 i_3272 (.ZN (n_2369), .A (n_68), .B1 (n_2274), .B2 (n_58));
OR2_X1 i_3271 (.ZN (n_2368), .A1 (n_58), .A2 (n_1132));
OAI22_X1 i_3270 (.ZN (n_2367), .A1 (n_2370), .A2 (n_2369), .B1 (n_68), .B2 (n_2368));
NAND2_X1 i_3268 (.ZN (n_2366), .A1 (n_2371), .A2 (n_2367));
XNOR2_X1 i_3267 (.ZN (n_2365), .A (n_2403), .B (n_2402));
NOR2_X1 i_3266 (.ZN (n_2364), .A1 (n_2366), .A2 (n_2365));
OR2_X1 i_3265 (.ZN (n_2363), .A1 (n_10), .A2 (n_11));
NAND2_X1 i_3264 (.ZN (n_2362), .A1 (inputA[0]), .A2 (inputB[4]));
OAI21_X1 i_3263 (.ZN (n_2361), .A (n_2409), .B1 (n_2363), .B2 (n_2362));
NAND2_X1 i_3262 (.ZN (n_2360), .A1 (n_2369), .A2 (n_2361));
OAI21_X1 i_3261 (.ZN (n_2359), .A (n_2360), .B1 (n_2369), .B2 (n_2361));
NAND2_X1 i_3260 (.ZN (n_2358), .A1 (inputA[3]), .A2 (inputB[2]));
XNOR2_X1 i_3259 (.ZN (n_2357), .A (n_2406), .B (n_2358));
OAI21_X1 i_3258 (.ZN (n_2356), .A (n_2360), .B1 (n_2359), .B2 (n_2357));
NAND2_X1 i_3257 (.ZN (n_2355), .A1 (n_2364), .A2 (n_2356));
INV_X1 i_3256 (.ZN (n_2354), .A (n_2355));
NAND2_X1 i_3255 (.ZN (n_2353), .A1 (inputA[3]), .A2 (inputB[4]));
XOR2_X1 i_3254 (.Z (n_2352), .A (n_2284), .B (n_2353));
XOR2_X1 i_3253 (.Z (n_2351), .A (n_2279), .B (n_2280));
XOR2_X1 i_3252 (.Z (n_2350), .A (n_2352), .B (n_2351));
AOI22_X1 i_3251 (.ZN (n_2349), .A1 (n_2352), .A2 (n_2351), .B1 (n_2354), .B2 (n_2350));
NAND2_X1 i_3250 (.ZN (n_2348), .A1 (inputA[2]), .A2 (inputB[6]));
XNOR2_X1 i_3249 (.ZN (n_2347), .A (n_2242), .B (n_2348));
NAND2_X1 i_3248 (.ZN (n_2346), .A1 (inputA[0]), .A2 (inputB[8]));
XOR2_X1 i_3247 (.Z (n_2345), .A (n_2347), .B (n_2346));
XOR2_X1 i_3246 (.Z (n_2344), .A (n_2228), .B (n_2227));
NOR2_X1 i_3245 (.ZN (n_2343), .A1 (n_2345), .A2 (n_2344));
AOI21_X1 i_3244 (.ZN (n_2342), .A (n_2343), .B1 (n_2345), .B2 (n_2344));
INV_X1 i_3243 (.ZN (n_2341), .A (n_2342));
XOR2_X1 i_3242 (.Z (n_2340), .A (n_2218), .B (n_2217));
NOR2_X1 i_3241 (.ZN (n_2339), .A1 (n_2341), .A2 (n_2340));
AOI21_X1 i_3240 (.ZN (n_2338), .A (n_2339), .B1 (n_2341), .B2 (n_2340));
NOR2_X1 i_3239 (.ZN (n_2337), .A1 (n_2349), .A2 (n_2338));
NAND2_X1 i_3238 (.ZN (n_2336), .A1 (n_2372), .A2 (n_2337));
INV_X1 i_3237 (.ZN (n_2335), .A (n_2336));
XNOR2_X1 i_3236 (.ZN (n_2331), .A (n_2262), .B (n_2261));
NAND2_X1 i_3235 (.ZN (n_2330), .A1 (inputA[6]), .A2 (inputB[3]));
XOR2_X1 i_3234 (.Z (n_2329), .A (n_2257), .B (n_2330));
OAI22_X1 i_3233 (.ZN (n_2328), .A1 (n_2242), .A2 (n_2348), .B1 (n_2347), .B2 (n_2346));
XOR2_X1 i_3232 (.Z (n_2327), .A (n_2329), .B (n_2328));
NAND2_X1 i_3231 (.ZN (n_2326), .A1 (inputA[3]), .A2 (inputB[6]));
XOR2_X1 i_3230 (.Z (n_2325), .A (n_2243), .B (n_2326));
NOR2_X1 i_3229 (.ZN (n_2324), .A1 (n_2343), .A2 (n_2339));
XOR2_X1 i_3228 (.Z (n_2323), .A (n_2327), .B (n_2325));
NOR2_X1 i_3227 (.ZN (n_2322), .A1 (n_2324), .A2 (n_2323));
AOI21_X1 i_3226 (.ZN (n_2321), .A (n_2322), .B1 (n_2324), .B2 (n_2323));
AOI21_X1 i_3225 (.ZN (n_2320), .A (n_2322), .B1 (n_2331), .B2 (n_2321));
NAND2_X1 i_3224 (.ZN (n_2319), .A1 (n_2335), .A2 (n_2320));
INV_X1 i_3223 (.ZN (n_2318), .A (n_2232));
NAND2_X1 i_3222 (.ZN (n_2317), .A1 (inputB[3]), .A2 (inputA[7]));
NAND2_X1 i_3221 (.ZN (n_2316), .A1 (inputB[2]), .A2 (inputA[8]));
XOR2_X1 i_3220 (.Z (n_2315), .A (n_2317), .B (n_2316));
INV_X1 i_3219 (.ZN (n_2314), .A (n_2315));
NAND2_X1 i_3218 (.ZN (n_2313), .A1 (inputB[4]), .A2 (inputA[6]));
XNOR2_X1 i_3217 (.ZN (n_2312), .A (n_2315), .B (n_2313));
XOR2_X1 i_3216 (.Z (n_2292), .A (n_2252), .B (n_2255));
XOR2_X1 i_3215 (.Z (n_2291), .A (n_2312), .B (n_2292));
NAND2_X1 i_3214 (.ZN (n_2290), .A1 (inputB[5]), .A2 (inputA[5]));
XNOR2_X1 i_3213 (.ZN (n_2289), .A (n_2203), .B (n_2290));
NAND2_X1 i_3212 (.ZN (n_2288), .A1 (inputB[7]), .A2 (inputA[3]));
XOR2_X1 i_3211 (.Z (n_2287), .A (n_2289), .B (n_2288));
XNOR2_X1 i_3210 (.ZN (n_2286), .A (n_2291), .B (n_2287));
NAND2_X1 i_3209 (.ZN (n_2285), .A1 (inputB[2]), .A2 (inputA[5]));
XNOR2_X1 i_3208 (.ZN (n_2284), .A (n_2221), .B (n_2285));
NAND2_X1 i_3207 (.ZN (n_2283), .A1 (inputB[6]), .A2 (inputA[0]));
AOI22_X1 i_3206 (.ZN (n_2282), .A1 (inputB[6]), .A2 (inputA[1]), .B1 (inputB[7]), .B2 (inputA[0]));
INV_X1 i_3205 (.ZN (n_2281), .A (n_2282));
OAI21_X1 i_3204 (.ZN (n_2280), .A (n_2281), .B1 (n_2242), .B2 (n_2283));
NAND2_X1 i_3203 (.ZN (n_2279), .A1 (inputB[5]), .A2 (inputA[2]));
OAI22_X1 i_3202 (.ZN (n_2278), .A1 (n_2242), .A2 (n_2283), .B1 (n_2280), .B2 (n_2279));
OAI33_X1 i_3201 (.ZN (n_2277), .A1 (n_1724), .A2 (n_690), .A3 (n_2284), .B1 (n_685)
    , .B2 (n_1132), .B3 (n_2285));
NOR2_X1 i_3200 (.ZN (n_2276), .A1 (n_2278), .A2 (n_2277));
AOI21_X1 i_3199 (.ZN (n_2275), .A (n_2276), .B1 (n_2278), .B2 (n_2277));
NAND2_X1 i_3198 (.ZN (n_2274), .A1 (inputB[1]), .A2 (inputA[4]));
NOR2_X1 i_3197 (.ZN (n_2273), .A1 (n_2285), .A2 (n_2274));
AOI22_X1 i_3196 (.ZN (n_2272), .A1 (inputB[1]), .A2 (inputA[5]), .B1 (inputB[2]), .B2 (inputA[4]));
NOR2_X1 i_3195 (.ZN (n_2271), .A1 (n_2273), .A2 (n_2272));
NOR2_X1 i_3194 (.ZN (n_2270), .A1 (n_1724), .A2 (n_685));
AOI21_X1 i_3193 (.ZN (n_2269), .A (n_2273), .B1 (n_2271), .B2 (n_2270));
INV_X1 i_3192 (.ZN (n_2268), .A (n_2269));
NOR2_X1 i_3191 (.ZN (n_2267), .A1 (n_63), .A2 (n_1349));
XOR2_X1 i_3190 (.Z (n_2266), .A (n_2318), .B (n_2267));
AOI22_X1 i_3189 (.ZN (n_2265), .A1 (n_2318), .A2 (n_2267), .B1 (n_2268), .B2 (n_2266));
AOI21_X1 i_3188 (.ZN (n_2264), .A (n_2276), .B1 (n_2275), .B2 (n_2265));
XOR2_X1 i_3187 (.Z (n_2263), .A (n_2238), .B (n_2237));
XOR2_X1 i_3186 (.Z (n_2262), .A (n_2264), .B (n_2263));
AOI21_X1 i_3185 (.ZN (n_2261), .A (n_2215), .B1 (n_2222), .B2 (n_2216));
AOI22_X1 i_3184 (.ZN (n_2260), .A1 (n_2264), .A2 (n_2263), .B1 (n_2262), .B2 (n_2261));
XOR2_X1 i_3183 (.Z (n_2259), .A (n_2286), .B (n_2260));
NAND2_X1 i_3182 (.ZN (n_2258), .A1 (inputB[2]), .A2 (inputA[7]));
XNOR2_X1 i_3181 (.ZN (n_2257), .A (n_2231), .B (n_2258));
OAI33_X1 i_3180 (.ZN (n_2255), .A1 (n_685), .A2 (n_1349), .A3 (n_2257), .B1 (n_2231)
    , .B2 (n_1219), .B3 (n_864));
OR2_X1 i_3179 (.ZN (n_2254), .A1 (n_63), .A2 (n_1894));
NOR2_X1 i_3178 (.ZN (n_2253), .A1 (n_2181), .A2 (n_2254));
AOI21_X1 i_3177 (.ZN (n_2252), .A (n_2253), .B1 (n_2181), .B2 (n_2254));
AOI21_X1 i_3176 (.ZN (n_2251), .A (n_2253), .B1 (n_2255), .B2 (n_2252));
XNOR2_X1 i_3175 (.ZN (n_2250), .A (n_2176), .B (n_2175));
NOR2_X1 i_3174 (.ZN (n_2249), .A1 (n_2251), .A2 (n_2250));
AOI21_X1 i_3173 (.ZN (n_2248), .A (n_2249), .B1 (n_2251), .B2 (n_2250));
XOR2_X1 i_3172 (.Z (n_2247), .A (n_2184), .B (n_2183));
XOR2_X1 i_3171 (.Z (n_2246), .A (n_2248), .B (n_2247));
NAND2_X1 i_3170 (.ZN (n_2245), .A1 (inputB[4]), .A2 (inputA[5]));
NAND2_X1 i_3169 (.ZN (n_2244), .A1 (inputB[5]), .A2 (inputA[4]));
XNOR2_X1 i_3168 (.ZN (n_2243), .A (n_2245), .B (n_2244));
NAND2_X1 i_3167 (.ZN (n_2242), .A1 (inputB[7]), .A2 (inputA[1]));
NAND2_X1 i_3166 (.ZN (n_2241), .A1 (inputB[8]), .A2 (inputA[2]));
AOI22_X1 i_3165 (.ZN (n_2240), .A1 (inputB[7]), .A2 (inputA[2]), .B1 (inputB[8]), .B2 (inputA[1]));
INV_X1 i_3164 (.ZN (n_2239), .A (n_2240));
OAI21_X1 i_3163 (.ZN (n_2238), .A (n_2239), .B1 (n_2242), .B2 (n_2241));
NAND2_X1 i_3162 (.ZN (n_2237), .A1 (inputB[9]), .A2 (inputA[0]));
OAI33_X1 i_3160 (.ZN (n_2236), .A1 (n_1724), .A2 (n_878), .A3 (n_2243), .B1 (n_1132)
    , .B2 (n_668), .B3 (n_2245));
OAI22_X1 i_3159 (.ZN (n_2235), .A1 (n_2242), .A2 (n_2241), .B1 (n_2238), .B2 (n_2237));
NAND2_X1 i_3158 (.ZN (n_2234), .A1 (n_2236), .A2 (n_2235));
OAI21_X1 i_3157 (.ZN (n_2233), .A (n_2234), .B1 (n_2236), .B2 (n_2235));
NAND2_X1 i_3156 (.ZN (n_2232), .A1 (inputB[0]), .A2 (inputA[7]));
NAND2_X1 i_3155 (.ZN (n_2231), .A1 (inputB[1]), .A2 (inputA[8]));
NOR2_X1 i_3154 (.ZN (n_2230), .A1 (n_2232), .A2 (n_2231));
AOI22_X1 i_3153 (.ZN (n_2229), .A1 (inputB[1]), .A2 (inputA[7]), .B1 (inputB[0]), .B2 (inputA[8]));
NOR2_X1 i_3152 (.ZN (n_2228), .A1 (n_2230), .A2 (n_2229));
NOR2_X1 i_3151 (.ZN (n_2227), .A1 (n_1219), .A2 (n_1349));
OR2_X1 i_3150 (.ZN (n_2226), .A1 (n_62), .A2 (n_1894));
AOI21_X1 i_3149 (.ZN (n_2225), .A (n_2230), .B1 (n_2228), .B2 (n_2227));
NOR2_X1 i_3148 (.ZN (n_2224), .A1 (n_2226), .A2 (n_2225));
AOI21_X1 i_3147 (.ZN (n_2223), .A (n_2224), .B1 (n_2226), .B2 (n_2225));
INV_X1 i_3146 (.ZN (n_2222), .A (n_2223));
NAND2_X1 i_3145 (.ZN (n_2221), .A1 (inputB[3]), .A2 (inputA[4]));
NOR2_X1 i_3144 (.ZN (n_2220), .A1 (n_2245), .A2 (n_2221));
AOI22_X1 i_3143 (.ZN (n_2219), .A1 (inputB[3]), .A2 (inputA[5]), .B1 (inputB[4]), .B2 (inputA[4]));
NOR2_X1 i_3142 (.ZN (n_2218), .A1 (n_2220), .A2 (n_2219));
NOR2_X1 i_3141 (.ZN (n_2217), .A1 (n_1724), .A2 (n_668));
AOI21_X1 i_3140 (.ZN (n_2216), .A (n_2220), .B1 (n_2218), .B2 (n_2217));
NOR2_X1 i_3139 (.ZN (n_2215), .A1 (n_2222), .A2 (n_2216));
NOR2_X1 i_3138 (.ZN (n_2214), .A1 (n_2224), .A2 (n_2215));
OAI21_X1 i_3137 (.ZN (n_2208), .A (n_2234), .B1 (n_2233), .B2 (n_2214));
XOR2_X1 i_3136 (.Z (n_2207), .A (n_2199), .B (n_2198));
XNOR2_X1 i_3135 (.ZN (n_2206), .A (n_2190), .B (n_2189));
XOR2_X1 i_3134 (.Z (n_2205), .A (n_2207), .B (n_2206));
XOR2_X1 i_3133 (.Z (n_2204), .A (n_2208), .B (n_2205));
NAND2_X1 i_3132 (.ZN (n_2203), .A1 (inputA[4]), .A2 (inputB[6]));
NAND2_X1 i_3131 (.ZN (n_2202), .A1 (inputA[5]), .A2 (inputB[7]));
NOR2_X1 i_3130 (.ZN (n_2201), .A1 (n_2203), .A2 (n_2202));
AOI22_X1 i_3129 (.ZN (n_2200), .A1 (inputA[4]), .A2 (inputB[7]), .B1 (inputA[5]), .B2 (inputB[6]));
NOR2_X1 i_3128 (.ZN (n_2199), .A1 (n_2201), .A2 (n_2200));
NOR2_X1 i_3127 (.ZN (n_2198), .A1 (n_1724), .A2 (n_669));
AOI21_X1 i_3126 (.ZN (n_2197), .A (n_2201), .B1 (n_2199), .B2 (n_2198));
INV_X1 i_3125 (.ZN (n_2196), .A (n_2197));
NAND2_X1 i_3124 (.ZN (n_2195), .A1 (inputA[1]), .A2 (inputB[9]));
NAND2_X1 i_3123 (.ZN (n_2194), .A1 (inputA[2]), .A2 (inputB[10]));
NOR2_X1 i_3122 (.ZN (n_2193), .A1 (n_2195), .A2 (n_2194));
INV_X1 i_3121 (.ZN (n_2192), .A (n_2193));
AOI22_X1 i_3120 (.ZN (n_2191), .A1 (inputA[1]), .A2 (inputB[10]), .B1 (inputA[2]), .B2 (inputB[9]));
NOR2_X1 i_3119 (.ZN (n_2190), .A1 (n_2193), .A2 (n_2191));
NAND2_X1 i_3118 (.ZN (n_2189), .A1 (inputA[0]), .A2 (inputB[11]));
AOI21_X1 i_3117 (.ZN (n_2188), .A (n_2191), .B1 (n_2192), .B2 (n_2189));
XOR2_X1 i_3116 (.Z (n_2187), .A (n_2196), .B (n_2188));
NAND2_X1 i_3115 (.ZN (n_2186), .A1 (inputB[3]), .A2 (inputA[8]));
NAND2_X1 i_3114 (.ZN (n_2185), .A1 (inputB[4]), .A2 (inputA[7]));
XNOR2_X1 i_3113 (.ZN (n_2184), .A (n_2186), .B (n_2185));
NAND2_X1 i_3112 (.ZN (n_2183), .A1 (inputB[5]), .A2 (inputA[6]));
OAI22_X1 i_3111 (.ZN (n_2182), .A1 (n_2186), .A2 (n_2185), .B1 (n_2184), .B2 (n_2183));
NAND2_X1 i_3110 (.ZN (n_2181), .A1 (inputB[0]), .A2 (inputA[10]));
NAND2_X1 i_3109 (.ZN (n_2180), .A1 (inputB[1]), .A2 (inputA[11]));
NOR2_X1 i_3108 (.ZN (n_2179), .A1 (n_2181), .A2 (n_2180));
AOI22_X1 i_3107 (.ZN (n_2178), .A1 (inputB[1]), .A2 (inputA[10]), .B1 (inputB[0]), .B2 (inputA[11]));
NOR2_X1 i_3106 (.ZN (n_2176), .A1 (n_2179), .A2 (n_2178));
NOR2_X1 i_3105 (.ZN (n_2175), .A1 (n_1219), .A2 (n_1894));
AOI21_X1 i_3104 (.ZN (n_2174), .A (n_2179), .B1 (n_2176), .B2 (n_2175));
NOR2_X1 i_3103 (.ZN (n_2173), .A1 (n_62), .A2 (n_667));
XNOR2_X1 i_3102 (.ZN (n_2172), .A (n_2182), .B (n_2174));
NAND2_X1 i_3101 (.ZN (n_2171), .A1 (n_2173), .A2 (n_2172));
OAI21_X1 i_3100 (.ZN (n_2170), .A (n_2171), .B1 (n_2173), .B2 (n_2172));
INV_X1 i_3099 (.ZN (n_2169), .A (n_16));
INV_X1 i_3098 (.ZN (n_2168), .A (n_1858));
XOR2_X1 i_3097 (.Z (n_2167), .A (n_1829), .B (n_1828));
XNOR2_X1 i_3096 (.ZN (n_2166), .A (n_1840), .B (n_1839));
XOR2_X1 i_3095 (.Z (n_2165), .A (n_2167), .B (n_2166));
NAND2_X1 i_3094 (.ZN (n_2164), .A1 (n_2169), .A2 (n_1824));
OAI21_X1 i_3093 (.ZN (n_2163), .A (n_2164), .B1 (n_2169), .B2 (n_1824));
NAND2_X1 i_3092 (.ZN (n_2162), .A1 (inputA[0]), .A2 (inputB[15]));
XNOR2_X1 i_3091 (.ZN (n_2161), .A (n_2163), .B (n_2162));
AOI22_X1 i_3090 (.ZN (n_2149), .A1 (n_2167), .A2 (n_2166), .B1 (n_2165), .B2 (n_2161));
INV_X1 i_3089 (.ZN (n_2148), .A (n_2149));
XOR2_X1 i_3088 (.Z (n_2147), .A (n_1834), .B (n_1826));
NAND2_X1 i_3087 (.ZN (n_2146), .A1 (n_2148), .A2 (n_2147));
OAI21_X1 i_3086 (.ZN (n_2141), .A (n_2146), .B1 (n_2148), .B2 (n_2147));
NAND2_X1 i_3085 (.ZN (n_2140), .A1 (inputA[6]), .A2 (inputB[6]));
NOR2_X1 i_3084 (.ZN (n_2139), .A1 (n_1843), .A2 (n_2140));
AOI22_X1 i_3083 (.ZN (n_2138), .A1 (inputA[7]), .A2 (inputB[6]), .B1 (inputA[6]), .B2 (inputB[7]));
NOR2_X1 i_3082 (.ZN (n_2137), .A1 (n_2139), .A2 (n_2138));
NAND2_X1 i_3081 (.ZN (n_2136), .A1 (inputA[8]), .A2 (inputB[5]));
NAND2_X1 i_3080 (.ZN (n_2135), .A1 (inputA[10]), .A2 (inputB[2]));
NAND2_X1 i_3079 (.ZN (n_2134), .A1 (inputA[11]), .A2 (inputB[3]));
NOR2_X1 i_3078 (.ZN (n_2133), .A1 (n_2135), .A2 (n_2134));
AOI22_X1 i_3077 (.ZN (n_2132), .A1 (inputA[10]), .A2 (inputB[3]), .B1 (inputA[11]), .B2 (inputB[2]));
NOR2_X1 i_3076 (.ZN (n_2131), .A1 (n_2133), .A2 (n_2132));
NOR2_X1 i_3075 (.ZN (n_2130), .A1 (n_690), .A2 (n_1894));
OAI22_X1 i_3074 (.ZN (n_2129), .A1 (n_1843), .A2 (n_2140), .B1 (n_2138), .B2 (n_2136));
AOI21_X1 i_3073 (.ZN (n_2128), .A (n_2133), .B1 (n_2131), .B2 (n_2130));
INV_X1 i_3072 (.ZN (n_2127), .A (n_2128));
XOR2_X1 i_3071 (.Z (n_2126), .A (n_2129), .B (n_2127));
NAND2_X1 i_3070 (.ZN (n_2125), .A1 (inputA[4]), .A2 (inputB[9]));
NAND2_X1 i_3069 (.ZN (n_2124), .A1 (inputA[5]), .A2 (inputB[8]));
XNOR2_X1 i_3068 (.ZN (n_2122), .A (n_2125), .B (n_2124));
NAND2_X1 i_3067 (.ZN (n_2121), .A1 (inputA[3]), .A2 (inputB[10]));
OAI22_X1 i_3066 (.ZN (n_2120), .A1 (n_2125), .A2 (n_2124), .B1 (n_2122), .B2 (n_2121));
AOI22_X1 i_3065 (.ZN (n_2119), .A1 (n_2129), .A2 (n_2127), .B1 (n_2126), .B2 (n_2120));
NAND2_X1 i_3064 (.ZN (n_2118), .A1 (inputA[14]), .A2 (inputB[1]));
NAND2_X1 i_3063 (.ZN (n_2117), .A1 (inputA[13]), .A2 (inputB[2]));
XNOR2_X1 i_3062 (.ZN (n_2116), .A (n_2118), .B (n_2117));
NAND2_X1 i_3061 (.ZN (n_2115), .A1 (inputA[12]), .A2 (inputB[3]));
XOR2_X1 i_3060 (.Z (n_2114), .A (n_2116), .B (n_2115));
NAND2_X1 i_3059 (.ZN (n_2113), .A1 (inputA[9]), .A2 (inputB[6]));
XOR2_X1 i_3058 (.Z (n_2112), .A (n_1845), .B (n_2113));
NOR2_X1 i_3057 (.ZN (n_2111), .A1 (n_2114), .A2 (n_2112));
AOI21_X1 i_3056 (.ZN (n_2110), .A (n_2111), .B1 (n_2114), .B2 (n_2112));
AOI21_X1 i_3055 (.ZN (n_2109), .A (n_2111), .B1 (n_2119), .B2 (n_2110));
AOI21_X1 i_3054 (.ZN (n_2108), .A (n_2168), .B1 (n_1860), .B2 (n_1859));
OAI21_X1 i_3053 (.ZN (n_2107), .A (n_2146), .B1 (n_2141), .B2 (n_2109));
NAND2_X1 i_3052 (.ZN (n_2106), .A1 (n_2108), .A2 (n_2107));
OAI21_X1 i_3051 (.ZN (n_2105), .A (n_2106), .B1 (n_2108), .B2 (n_2107));
NAND2_X1 i_3050 (.ZN (n_2104), .A1 (inputA[15]), .A2 (inputB[0]));
OAI22_X1 i_3049 (.ZN (n_2103), .A1 (n_62), .A2 (n_865), .B1 (n_63), .B2 (n_478));
INV_X1 i_3048 (.ZN (n_2102), .A (n_2103));
OAI22_X1 i_3047 (.ZN (n_2101), .A1 (n_2118), .A2 (n_2117), .B1 (n_2116), .B2 (n_2115));
NOR2_X1 i_3046 (.ZN (n_2100), .A1 (n_1893), .A2 (n_2104));
OAI21_X1 i_3045 (.ZN (n_2099), .A (n_2103), .B1 (n_2101), .B2 (n_2100));
INV_X1 i_3044 (.ZN (n_2098), .A (n_2099));
XOR2_X1 i_3043 (.Z (n_2097), .A (n_1891), .B (n_1890));
XNOR2_X1 i_3042 (.ZN (n_2096), .A (n_2098), .B (n_2097));
XNOR2_X1 i_3041 (.ZN (n_2095), .A (n_1886), .B (n_1870));
NOR2_X1 i_3039 (.ZN (n_2094), .A1 (n_2096), .A2 (n_2095));
AOI21_X1 i_3038 (.ZN (n_2093), .A (n_2094), .B1 (n_2096), .B2 (n_2095));
OAI21_X1 i_3037 (.ZN (n_2092), .A (n_2106), .B1 (n_2105), .B2 (n_2093));
XNOR2_X1 i_3036 (.ZN (n_2091), .A (n_1864), .B (n_1857));
NOR2_X1 i_3035 (.ZN (n_2090), .A1 (n_2092), .A2 (n_2091));
AOI21_X1 i_3034 (.ZN (n_2083), .A (n_2090), .B1 (n_2092), .B2 (n_2091));
XOR2_X1 i_3033 (.Z (n_2082), .A (n_2015), .B (n_2014));
NAND2_X1 i_3032 (.ZN (n_2081), .A1 (n_1823), .A2 (n_1773));
OAI21_X1 i_3031 (.ZN (n_2080), .A (n_2081), .B1 (n_1823), .B2 (n_1773));
NAND2_X1 i_3030 (.ZN (n_2079), .A1 (inputA[0]), .A2 (inputB[17]));
OAI21_X1 i_3029 (.ZN (n_2078), .A (n_2081), .B1 (n_2080), .B2 (n_2079));
XOR2_X1 i_3028 (.Z (n_2077), .A (n_2082), .B (n_2078));
NOR2_X1 i_3027 (.ZN (n_2076), .A1 (n_1847), .A2 (n_1735));
AOI22_X1 i_3026 (.ZN (n_2075), .A1 (inputA[10]), .A2 (inputB[6]), .B1 (inputA[11]), .B2 (inputB[5]));
NOR2_X1 i_3025 (.ZN (n_2074), .A1 (n_2076), .A2 (n_2075));
NOR2_X1 i_3024 (.ZN (n_2073), .A1 (n_1894), .A2 (n_879));
AOI21_X1 i_3023 (.ZN (n_2072), .A (n_2076), .B1 (n_2074), .B2 (n_2073));
NOR2_X1 i_3022 (.ZN (n_2071), .A1 (n_1888), .A2 (n_2117));
AOI22_X1 i_3021 (.ZN (n_2070), .A1 (inputA[13]), .A2 (inputB[3]), .B1 (inputA[14]), .B2 (inputB[2]));
NOR2_X1 i_3020 (.ZN (n_2069), .A1 (n_2071), .A2 (n_2070));
NOR2_X1 i_3019 (.ZN (n_2068), .A1 (n_690), .A2 (n_667));
AOI21_X1 i_3018 (.ZN (n_2067), .A (n_2071), .B1 (n_2069), .B2 (n_2068));
XNOR2_X1 i_3017 (.ZN (n_2066), .A (n_2072), .B (n_2067));
NOR3_X1 i_3016 (.ZN (n_2065), .A1 (n_1731), .A2 (n_669), .A3 (n_864));
AOI22_X1 i_3015 (.ZN (n_2064), .A1 (inputA[7]), .A2 (inputB[9]), .B1 (inputA[8]), .B2 (inputB[8]));
OR2_X1 i_3014 (.ZN (n_2063), .A1 (n_2065), .A2 (n_2064));
OR2_X1 i_3013 (.ZN (n_2062), .A1 (n_1349), .A2 (n_1131));
NOR2_X1 i_3012 (.ZN (n_2061), .A1 (n_2063), .A2 (n_2062));
NOR2_X1 i_3011 (.ZN (n_2060), .A1 (n_2065), .A2 (n_2061));
OAI22_X1 i_3010 (.ZN (n_2059), .A1 (n_2072), .A2 (n_2067), .B1 (n_2066), .B2 (n_2060));
XOR2_X1 i_3009 (.Z (n_2058), .A (n_2077), .B (n_2059));
AOI21_X1 i_3008 (.ZN (n_2057), .A (n_2094), .B1 (n_2098), .B2 (n_2097));
XNOR2_X1 i_3007 (.ZN (n_2056), .A (n_2058), .B (n_2057));
AOI21_X1 i_3006 (.ZN (n_2055), .A (n_2061), .B1 (n_2063), .B2 (n_2062));
XOR2_X1 i_3005 (.Z (n_2054), .A (n_1813), .B (n_1812));
NOR2_X1 i_3004 (.ZN (n_2053), .A1 (n_2055), .A2 (n_2054));
AOI21_X1 i_3003 (.ZN (n_2052), .A (n_2053), .B1 (n_2055), .B2 (n_2054));
XNOR2_X1 i_3002 (.ZN (n_2051), .A (n_1821), .B (n_1820));
XOR2_X1 i_3001 (.Z (n_2050), .A (n_2066), .B (n_2060));
AOI21_X1 i_3000 (.ZN (n_2049), .A (n_2053), .B1 (n_2052), .B2 (n_2051));
NOR2_X1 i_2999 (.ZN (n_2048), .A1 (n_2050), .A2 (n_2049));
AOI21_X1 i_2998 (.ZN (n_2047), .A (n_2048), .B1 (n_2050), .B2 (n_2049));
NOR2_X1 i_2997 (.ZN (n_2046), .A1 (n_2102), .A2 (n_2100));
XNOR2_X1 i_2996 (.ZN (n_2045), .A (n_2101), .B (n_2046));
XNOR2_X1 i_2995 (.ZN (n_2044), .A (n_2069), .B (n_2068));
NOR2_X1 i_2994 (.ZN (n_2043), .A1 (n_2045), .A2 (n_2044));
AOI21_X1 i_2993 (.ZN (n_2042), .A (n_2043), .B1 (n_2045), .B2 (n_2044));
XOR2_X1 i_2992 (.Z (n_2041), .A (n_2074), .B (n_2073));
AOI21_X1 i_2991 (.ZN (n_2040), .A (n_2043), .B1 (n_2042), .B2 (n_2041));
AOI21_X1 i_2990 (.ZN (n_2039), .A (n_2048), .B1 (n_2047), .B2 (n_2040));
XOR2_X1 i_2989 (.Z (n_2038), .A (n_2056), .B (n_2039));
AOI21_X1 i_2988 (.ZN (n_2037), .A (n_2090), .B1 (n_2083), .B2 (n_2038));
INV_X1 i_2987 (.ZN (n_2036), .A (n_1917));
NOR2_X1 i_2986 (.ZN (n_2035), .A1 (n_1893), .A2 (n_1915));
AOI22_X1 i_2985 (.ZN (n_2016), .A1 (inputB[1]), .A2 (inputA[17]), .B1 (inputB[2]), .B2 (inputA[16]));
NOR2_X1 i_2984 (.ZN (n_2015), .A1 (n_2035), .A2 (n_2016));
NOR2_X1 i_2983 (.ZN (n_2014), .A1 (n_685), .A2 (n_478));
NAND2_X1 i_2982 (.ZN (n_2013), .A1 (inputB[1]), .A2 (inputA[19]));
NAND2_X1 i_2981 (.ZN (n_2012), .A1 (n_1889), .A2 (n_1869));
OAI21_X1 i_2980 (.ZN (n_2011), .A (n_2012), .B1 (n_1868), .B2 (n_1867));
AOI21_X1 i_2979 (.ZN (n_2010), .A (n_2035), .B1 (n_2015), .B2 (n_2014));
OAI22_X1 i_2978 (.ZN (n_2009), .A1 (n_63), .A2 (n_479), .B1 (n_62), .B2 (n_480));
OAI21_X1 i_2977 (.ZN (n_2008), .A (n_2009), .B1 (n_1867), .B2 (n_2013));
XOR2_X1 i_2976 (.Z (n_2007), .A (n_2010), .B (n_2008));
XOR2_X1 i_2975 (.Z (n_2006), .A (n_2011), .B (n_2007));
NOR2_X1 i_2974 (.ZN (n_2005), .A1 (n_1918), .A2 (n_2036));
XOR2_X1 i_2973 (.Z (n_2004), .A (n_1919), .B (n_2005));
AOI22_X1 i_2972 (.ZN (n_2003), .A1 (n_2011), .A2 (n_2007), .B1 (n_2006), .B2 (n_2004));
XOR2_X1 i_2971 (.Z (n_2002), .A (n_1926), .B (n_1927));
XNOR2_X1 i_2970 (.ZN (n_2001), .A (n_1911), .B (n_1912));
XOR2_X1 i_2969 (.Z (n_2000), .A (n_2002), .B (n_2001));
XNOR2_X1 i_2968 (.ZN (n_1999), .A (n_1899), .B (n_1900));
NAND2_X1 i_2967 (.ZN (n_1998), .A1 (n_2000), .A2 (n_1999));
OAI21_X1 i_2966 (.ZN (n_1995), .A (n_1998), .B1 (n_2002), .B2 (n_2001));
XOR2_X1 i_2965 (.Z (n_1994), .A (n_2003), .B (n_1995));
NAND2_X1 i_2964 (.ZN (n_1993), .A1 (inputB[4]), .A2 (inputA[14]));
XNOR2_X1 i_2963 (.ZN (n_1992), .A (n_1907), .B (n_1993));
NAND2_X1 i_2962 (.ZN (n_1991), .A1 (inputB[6]), .A2 (inputA[12]));
NOR2_X1 i_2961 (.ZN (n_1990), .A1 (n_1736), .A2 (n_1924));
AOI22_X1 i_2960 (.ZN (n_1989), .A1 (inputB[7]), .A2 (inputA[11]), .B1 (inputB[8]), .B2 (inputA[10]));
NOR2_X1 i_2959 (.ZN (n_1988), .A1 (n_1990), .A2 (n_1989));
NOR2_X1 i_2958 (.ZN (n_1987), .A1 (n_1894), .A2 (n_1127));
AOI21_X1 i_2957 (.ZN (n_1986), .A (n_1990), .B1 (n_1988), .B2 (n_1987));
INV_X1 i_2956 (.ZN (n_1985), .A (n_1986));
OAI22_X1 i_2955 (.ZN (n_1984), .A1 (n_1907), .A2 (n_1993), .B1 (n_1992), .B2 (n_1991));
XOR2_X1 i_2954 (.Z (n_1983), .A (n_1985), .B (n_1984));
NOR2_X1 i_2953 (.ZN (n_1982), .A1 (n_1732), .A2 (n_1897));
AOI22_X1 i_2952 (.ZN (n_1981), .A1 (inputB[10]), .A2 (inputA[8]), .B1 (inputB[11]), .B2 (inputA[7]));
NOR2_X1 i_2951 (.ZN (n_1980), .A1 (n_1982), .A2 (n_1981));
NOR2_X1 i_2950 (.ZN (n_1978), .A1 (n_1349), .A2 (n_880));
AOI21_X1 i_2949 (.ZN (n_1976), .A (n_1982), .B1 (n_1980), .B2 (n_1978));
INV_X1 i_2948 (.ZN (n_1975), .A (n_1976));
AOI22_X1 i_2947 (.ZN (n_1974), .A1 (n_1985), .A2 (n_1984), .B1 (n_1983), .B2 (n_1975));
OAI22_X1 i_2946 (.ZN (n_1973), .A1 (n_1867), .A2 (n_2013), .B1 (n_2010), .B2 (n_2008));
XNOR2_X1 i_2945 (.ZN (n_1972), .A (n_1974), .B (n_1973));
NAND2_X1 i_2944 (.ZN (n_1971), .A1 (inputB[0]), .A2 (inputA[20]));
XOR2_X1 i_2943 (.Z (n_1970), .A (n_2013), .B (n_1971));
INV_X1 i_2942 (.ZN (n_1969), .A (n_1970));
NAND2_X1 i_2941 (.ZN (n_1968), .A1 (inputB[2]), .A2 (inputA[18]));
XOR2_X1 i_2940 (.Z (n_1967), .A (n_1970), .B (n_1968));
XOR2_X1 i_2939 (.Z (n_1966), .A (n_1972), .B (n_1967));
XOR2_X1 i_2938 (.Z (n_1965), .A (n_1994), .B (n_1966));
NAND2_X1 i_2937 (.ZN (n_1964), .A1 (inputB[8]), .A2 (inputA[13]));
NOR2_X1 i_2936 (.ZN (n_1963), .A1 (n_1912), .A2 (n_1964));
AOI22_X1 i_2935 (.ZN (n_1962), .A1 (inputB[8]), .A2 (inputA[12]), .B1 (inputB[7]), .B2 (inputA[13]));
NOR2_X1 i_2934 (.ZN (n_1961), .A1 (n_1963), .A2 (n_1962));
XOR2_X1 i_2933 (.Z (n_1960), .A (n_1908), .B (n_1961));
NAND2_X1 i_2932 (.ZN (n_1948), .A1 (inputB[4]), .A2 (inputA[17]));
NOR2_X1 i_2931 (.ZN (n_1947), .A1 (n_1916), .A2 (n_1948));
AOI22_X1 i_2930 (.ZN (n_1946), .A1 (inputB[3]), .A2 (inputA[17]), .B1 (inputB[4]), .B2 (inputA[16]));
NOR2_X1 i_2929 (.ZN (n_1945), .A1 (n_1947), .A2 (n_1946));
NOR2_X1 i_2928 (.ZN (n_1944), .A1 (n_478), .A2 (n_668));
XNOR2_X1 i_2927 (.ZN (n_1940), .A (n_1945), .B (n_1944));
XOR2_X1 i_2926 (.Z (n_1939), .A (n_1960), .B (n_1940));
NAND2_X1 i_2925 (.ZN (n_1938), .A1 (inputB[10]), .A2 (inputA[11]));
NOR2_X1 i_2924 (.ZN (n_1937), .A1 (n_1925), .A2 (n_1938));
AOI22_X1 i_2923 (.ZN (n_1936), .A1 (inputB[9]), .A2 (inputA[11]), .B1 (inputB[10]), .B2 (inputA[10]));
NOR2_X1 i_2922 (.ZN (n_1935), .A1 (n_1937), .A2 (n_1936));
NAND2_X1 i_2921 (.ZN (n_1934), .A1 (inputB[11]), .A2 (inputA[9]));
XOR2_X1 i_2920 (.Z (n_1933), .A (n_1935), .B (n_1934));
XOR2_X1 i_2919 (.Z (n_1932), .A (n_1939), .B (n_1933));
XOR2_X1 i_2918 (.Z (n_1931), .A (n_1965), .B (n_1932));
XOR2_X1 i_2917 (.Z (n_1930), .A (n_1905), .B (n_1929));
XNOR2_X1 i_2916 (.ZN (n_1929), .A (n_1923), .B (n_1928));
OAI22_X1 i_2915 (.ZN (n_1928), .A1 (n_1926), .A2 (n_1927), .B1 (n_1924), .B2 (n_1925));
NAND2_X1 i_2914 (.ZN (n_1927), .A1 (inputA[9]), .A2 (inputB[10]));
XNOR2_X1 i_2913 (.ZN (n_1926), .A (n_1924), .B (n_1925));
NAND2_X1 i_2912 (.ZN (n_1925), .A1 (inputA[10]), .A2 (inputB[9]));
NAND2_X1 i_2911 (.ZN (n_1924), .A1 (inputA[11]), .A2 (inputB[8]));
XOR2_X1 i_2910 (.Z (n_1923), .A (n_1914), .B (n_1922));
OAI21_X1 i_2909 (.ZN (n_1922), .A (n_1917), .B1 (n_1918), .B2 (n_1919));
NOR2_X1 i_2908 (.ZN (n_1919), .A1 (n_690), .A2 (n_478));
NOR2_X1 i_2907 (.ZN (n_1918), .A1 (n_1915), .A2 (n_1916));
NAND2_X1 i_2905 (.ZN (n_1917), .A1 (n_1915), .A2 (n_1916));
NAND2_X1 i_2903 (.ZN (n_1916), .A1 (inputA[16]), .A2 (inputB[3]));
NAND2_X1 i_2902 (.ZN (n_1915), .A1 (inputA[17]), .A2 (inputB[2]));
AOI21_X1 i_2901 (.ZN (n_1914), .A (n_1909), .B1 (n_1911), .B2 (n_1913));
INV_X1 i_2900 (.ZN (n_1913), .A (n_1912));
NAND2_X1 i_2899 (.ZN (n_1912), .A1 (inputA[12]), .A2 (inputB[7]));
NOR2_X1 i_2897 (.ZN (n_1911), .A1 (n_1909), .A2 (n_1910));
AOI22_X1 i_2896 (.ZN (n_1910), .A1 (inputA[14]), .A2 (inputB[5]), .B1 (inputA[13]), .B2 (inputB[6]));
NOR2_X1 i_2895 (.ZN (n_1909), .A1 (n_1907), .A2 (n_1908));
NAND2_X1 i_2894 (.ZN (n_1908), .A1 (inputA[14]), .A2 (inputB[6]));
NAND2_X1 i_2893 (.ZN (n_1907), .A1 (inputB[5]), .A2 (inputA[13]));
XOR2_X1 i_2892 (.Z (n_1905), .A (n_1904), .B (n_1895));
XNOR2_X1 i_2891 (.ZN (n_1904), .A (n_1902), .B (n_1903));
AOI21_X1 i_2890 (.ZN (n_1903), .A (n_1789), .B1 (n_1791), .B2 (n_1725));
XOR2_X1 i_2889 (.Z (n_1902), .A (n_1901), .B (n_1896));
OAI22_X1 i_2888 (.ZN (n_1901), .A1 (n_1899), .A2 (n_1900), .B1 (n_1897), .B2 (n_1898));
NAND2_X1 i_2887 (.ZN (n_1900), .A1 (inputA[6]), .A2 (inputB[13]));
XNOR2_X1 i_2886 (.ZN (n_1899), .A (n_1897), .B (n_1898));
NAND2_X1 i_2885 (.ZN (n_1898), .A1 (inputA[7]), .A2 (inputB[12]));
NAND2_X1 i_2884 (.ZN (n_1897), .A1 (inputA[8]), .A2 (inputB[11]));
AOI21_X1 i_2883 (.ZN (n_1896), .A (n_1728), .B1 (n_1730), .B2 (n_1726));
AOI22_X1 i_2882 (.ZN (n_1895), .A1 (n_1785), .A2 (n_1782), .B1 (n_1772), .B2 (n_1786));
INV_X1 i_2881 (.ZN (n_1894), .A (inputA[9]));
NAND2_X1 i_2880 (.ZN (n_1893), .A1 (inputB[1]), .A2 (inputA[16]));
NAND2_X1 i_2879 (.ZN (n_1892), .A1 (inputB[0]), .A2 (inputA[17]));
XNOR2_X1 i_2878 (.ZN (n_1891), .A (n_1893), .B (n_1892));
NAND2_X1 i_2877 (.ZN (n_1890), .A1 (inputB[2]), .A2 (inputA[15]));
OAI22_X1 i_2876 (.ZN (n_1889), .A1 (n_1893), .A2 (n_1892), .B1 (n_1891), .B2 (n_1890));
NAND2_X1 i_2875 (.ZN (n_1888), .A1 (inputB[3]), .A2 (inputA[14]));
NAND2_X1 i_2874 (.ZN (n_1887), .A1 (inputB[4]), .A2 (inputA[13]));
XNOR2_X1 i_2873 (.ZN (n_1886), .A (n_1888), .B (n_1887));
NAND2_X1 i_2872 (.ZN (n_1870), .A1 (inputB[5]), .A2 (inputA[12]));
OAI22_X1 i_2871 (.ZN (n_1869), .A1 (n_1888), .A2 (n_1887), .B1 (n_1886), .B2 (n_1870));
XNOR2_X1 i_2870 (.ZN (n_1868), .A (n_1889), .B (n_1869));
NAND2_X1 i_2869 (.ZN (n_1867), .A1 (inputB[0]), .A2 (inputA[18]));
XOR2_X1 i_2868 (.Z (n_1866), .A (n_1764), .B (n_1771));
XOR2_X1 i_2867 (.Z (n_1865), .A (n_1868), .B (n_1867));
XNOR2_X1 i_2866 (.ZN (n_1864), .A (n_1866), .B (n_1865));
NAND2_X1 i_2865 (.ZN (n_1863), .A1 (inputB[11]), .A2 (inputA[6]));
XOR2_X1 i_2864 (.Z (n_1862), .A (n_1733), .B (n_1863));
XOR2_X1 i_2863 (.Z (n_1861), .A (n_1737), .B (n_1738));
XNOR2_X1 i_2862 (.ZN (n_1860), .A (n_1862), .B (n_1861));
XOR2_X1 i_2861 (.Z (n_1859), .A (n_1769), .B (n_1770));
OR2_X1 i_2860 (.ZN (n_1858), .A1 (n_1860), .A2 (n_1859));
OAI21_X1 i_2859 (.ZN (n_1857), .A (n_1858), .B1 (n_1862), .B2 (n_1861));
INV_X1 i_2858 (.ZN (n_1856), .A (n_1857));
NAND2_X1 i_2857 (.ZN (n_1847), .A1 (inputB[5]), .A2 (inputA[10]));
NAND2_X1 i_2856 (.ZN (n_1846), .A1 (inputB[4]), .A2 (inputA[11]));
XNOR2_X1 i_2855 (.ZN (n_1845), .A (n_1847), .B (n_1846));
NAND2_X1 i_2854 (.ZN (n_1844), .A1 (inputB[4]), .A2 (inputA[10]));
NAND2_X1 i_2853 (.ZN (n_1843), .A1 (inputB[7]), .A2 (inputA[7]));
NOR3_X1 i_2852 (.ZN (n_1842), .A1 (n_669), .A2 (n_1843), .A3 (n_1551));
AOI22_X1 i_2851 (.ZN (n_1841), .A1 (inputB[8]), .A2 (inputA[7]), .B1 (inputB[7]), .B2 (inputA[8]));
NOR2_X1 i_2850 (.ZN (n_1840), .A1 (n_1842), .A2 (n_1841));
NOR2_X1 i_2849 (.ZN (n_1839), .A1 (n_1349), .A2 (n_1127));
OAI33_X1 i_2848 (.ZN (n_1838), .A1 (n_1894), .A2 (n_878), .A3 (n_1845), .B1 (n_668)
    , .B2 (n_1136), .B3 (n_1844));
INV_X1 i_2847 (.ZN (n_1837), .A (n_1838));
AOI21_X1 i_2846 (.ZN (n_1836), .A (n_1842), .B1 (n_1840), .B2 (n_1839));
NOR2_X1 i_2845 (.ZN (n_1835), .A1 (n_1837), .A2 (n_1836));
AOI21_X1 i_2844 (.ZN (n_1834), .A (n_1835), .B1 (n_1837), .B2 (n_1836));
NAND2_X1 i_2843 (.ZN (n_1833), .A1 (inputB[11]), .A2 (inputA[3]));
NOR2_X1 i_2842 (.ZN (n_1832), .A1 (n_1765), .A2 (n_1833));
AOI22_X1 i_2841 (.ZN (n_1831), .A1 (inputB[11]), .A2 (inputA[4]), .B1 (inputB[12]), .B2 (inputA[3]));
NOR2_X1 i_2840 (.ZN (n_1829), .A1 (n_1832), .A2 (n_1831));
NAND2_X1 i_2839 (.ZN (n_1828), .A1 (inputB[10]), .A2 (inputA[5]));
OAI22_X1 i_2838 (.ZN (n_1827), .A1 (n_1765), .A2 (n_1833), .B1 (n_1831), .B2 (n_1828));
INV_X1 i_2837 (.ZN (n_1826), .A (n_1827));
AOI21_X1 i_2836 (.ZN (n_1825), .A (n_1835), .B1 (n_1834), .B2 (n_1827));
NOR2_X1 i_2835 (.ZN (n_1824), .A1 (n_1547), .A2 (n_586));
NOR2_X1 i_2834 (.ZN (n_1823), .A1 (n_67), .A2 (n_587));
AOI22_X1 i_2833 (.ZN (n_1822), .A1 (inputB[15]), .A2 (inputA[1]), .B1 (inputB[14]), .B2 (inputA[2]));
AOI21_X1 i_2832 (.ZN (n_1821), .A (n_1822), .B1 (n_1824), .B2 (n_1823));
NOR2_X1 i_2831 (.ZN (n_1820), .A1 (n_66), .A2 (n_588));
NAND2_X1 i_2830 (.ZN (n_1819), .A1 (inputB[11]), .A2 (inputA[5]));
XNOR2_X1 i_2829 (.ZN (n_1813), .A (n_1765), .B (n_1819));
NAND2_X1 i_2828 (.ZN (n_1812), .A1 (inputB[13]), .A2 (inputA[3]));
AOI22_X1 i_2827 (.ZN (n_1811), .A1 (n_1824), .A2 (n_1823), .B1 (n_1821), .B2 (n_1820));
INV_X1 i_2826 (.ZN (n_1810), .A (n_1811));
OAI22_X1 i_2825 (.ZN (n_1809), .A1 (n_1765), .A2 (n_1819), .B1 (n_1813), .B2 (n_1812));
NAND2_X1 i_2824 (.ZN (n_1808), .A1 (n_1810), .A2 (n_1809));
OAI21_X1 i_2823 (.ZN (n_1807), .A (n_1808), .B1 (n_1810), .B2 (n_1809));
OAI21_X1 i_2822 (.ZN (n_1806), .A (n_1808), .B1 (n_1825), .B2 (n_1807));
NAND2_X1 i_2821 (.ZN (n_1805), .A1 (inputB[15]), .A2 (inputA[3]));
XNOR2_X1 i_2820 (.ZN (n_1804), .A (n_1784), .B (n_1805));
OAI21_X1 i_2819 (.ZN (n_1803), .A (n_1781), .B1 (n_1780), .B2 (n_1727));
NAND2_X1 i_2818 (.ZN (n_1802), .A1 (n_1804), .A2 (n_1803));
OAI21_X1 i_2817 (.ZN (n_1801), .A (n_1802), .B1 (n_1804), .B2 (n_1803));
OAI22_X1 i_2816 (.ZN (n_1800), .A1 (n_1866), .A2 (n_1865), .B1 (n_1864), .B2 (n_1856));
OAI21_X1 i_2815 (.ZN (n_1799), .A (n_1802), .B1 (n_1806), .B2 (n_1801));
NAND2_X1 i_2814 (.ZN (n_1798), .A1 (n_1800), .A2 (n_1799));
OAI21_X1 i_2813 (.ZN (n_1797), .A (n_1798), .B1 (n_1800), .B2 (n_1799));
XOR2_X1 i_2812 (.Z (n_1796), .A (n_1787), .B (n_1793));
OAI21_X1 i_2811 (.ZN (n_1795), .A (n_1798), .B1 (n_1797), .B2 (n_1796));
AOI22_X1 i_2810 (.ZN (n_1794), .A1 (n_1787), .A2 (n_1793), .B1 (n_1788), .B2 (n_1792));
XOR2_X1 i_2809 (.Z (n_1793), .A (n_1788), .B (n_1792));
XOR2_X1 i_2808 (.Z (n_1792), .A (n_1791), .B (n_1725));
NOR2_X1 i_2807 (.ZN (n_1791), .A1 (n_1789), .A2 (n_1790));
AOI22_X1 i_2806 (.ZN (n_1790), .A1 (inputB[15]), .A2 (inputA[4]), .B1 (inputB[14]), .B2 (inputA[5]));
NOR2_X1 i_2805 (.ZN (n_1789), .A1 (n_1783), .A2 (n_1723));
XOR2_X1 i_2804 (.Z (n_1788), .A (n_1730), .B (n_1726));
XOR2_X1 i_2803 (.Z (n_1787), .A (n_1772), .B (n_1786));
XOR2_X1 i_2802 (.Z (n_1786), .A (n_1782), .B (n_1785));
OAI33_X1 i_2801 (.ZN (n_1785), .A1 (n_1784), .A2 (n_1724), .A3 (n_587), .B1 (n_859)
    , .B2 (n_671), .B3 (n_1783));
XNOR2_X1 i_2800 (.ZN (n_1784), .A (n_1783), .B (n_1766));
NAND2_X1 i_2799 (.ZN (n_1783), .A1 (inputB[14]), .A2 (inputA[4]));
NAND2_X1 i_2798 (.ZN (n_1782), .A1 (n_1781), .A2 (n_1777));
NAND2_X1 i_2797 (.ZN (n_1781), .A1 (n_1780), .A2 (n_1727));
NOR2_X1 i_2796 (.ZN (n_1780), .A1 (n_1778), .A2 (n_1779));
AOI22_X1 i_2795 (.ZN (n_1779), .A1 (inputA[1]), .A2 (inputB[17]), .B1 (inputA[2]), .B2 (inputB[16]));
INV_X1 i_2794 (.ZN (n_1778), .A (n_1777));
NAND2_X1 i_2793 (.ZN (n_1777), .A1 (n_1726), .A2 (n_1773));
NOR2_X1 i_2792 (.ZN (n_1773), .A1 (n_1547), .A2 (n_588));
OAI21_X1 i_2791 (.ZN (n_1772), .A (n_1763), .B1 (n_1764), .B2 (n_1771));
AOI21_X1 i_2790 (.ZN (n_1771), .A (n_1767), .B1 (n_1769), .B2 (n_1770));
NOR2_X1 i_2789 (.ZN (n_1770), .A1 (n_1724), .A2 (n_586));
NOR2_X1 i_2788 (.ZN (n_1769), .A1 (n_1767), .A2 (n_1768));
AOI22_X1 i_2787 (.ZN (n_1768), .A1 (inputA[4]), .A2 (inputB[13]), .B1 (inputA[5]), .B2 (inputB[12]));
NOR2_X1 i_2786 (.ZN (n_1767), .A1 (n_1765), .A2 (n_1766));
NAND2_X1 i_2785 (.ZN (n_1766), .A1 (inputB[13]), .A2 (inputA[5]));
NAND2_X1 i_2784 (.ZN (n_1765), .A1 (inputA[4]), .A2 (inputB[12]));
OAI21_X1 i_2783 (.ZN (n_1764), .A (n_1763), .B1 (n_1739), .B2 (n_1740));
NAND2_X1 i_2782 (.ZN (n_1763), .A1 (n_1739), .A2 (n_1740));
OAI22_X1 i_2781 (.ZN (n_1740), .A1 (n_1737), .A2 (n_1738), .B1 (n_1735), .B2 (n_1736));
OAI33_X1 i_2780 (.ZN (n_1739), .A1 (n_1733), .A2 (n_1349), .A3 (n_670), .B1 (n_1551)
    , .B2 (n_1127), .B3 (n_1732));
NAND2_X1 i_2779 (.ZN (n_1738), .A1 (inputA[9]), .A2 (inputB[8]));
XNOR2_X1 i_2778 (.ZN (n_1737), .A (n_1735), .B (n_1736));
NAND2_X1 i_2777 (.ZN (n_1736), .A1 (inputA[10]), .A2 (inputB[7]));
NAND2_X1 i_2776 (.ZN (n_1735), .A1 (inputA[11]), .A2 (inputB[6]));
XNOR2_X1 i_2775 (.ZN (n_1733), .A (n_1731), .B (n_1732));
NAND2_X1 i_2774 (.ZN (n_1732), .A1 (inputA[7]), .A2 (inputB[10]));
NAND2_X1 i_2773 (.ZN (n_1731), .A1 (inputA[8]), .A2 (inputB[9]));
NOR2_X1 i_2772 (.ZN (n_1730), .A1 (n_1728), .A2 (n_1729));
AOI22_X1 i_2771 (.ZN (n_1729), .A1 (inputB[18]), .A2 (inputA[1]), .B1 (inputA[0]), .B2 (inputB[19]));
AND3_X1 i_2770 (.ZN (n_1728), .A1 (n_1727), .A2 (inputB[19]), .A3 (inputA[1]));
NOR2_X1 i_2769 (.ZN (n_1727), .A1 (n_66), .A2 (n_400));
NOR2_X1 i_2768 (.ZN (n_1726), .A1 (n_67), .A2 (n_881));
NOR2_X1 i_2767 (.ZN (n_1725), .A1 (n_1724), .A2 (n_588));
INV_X1 i_2766 (.ZN (n_1724), .A (inputA[3]));
NAND2_X1 i_2765 (.ZN (n_1723), .A1 (inputB[15]), .A2 (inputA[5]));
XOR2_X1 i_2764 (.Z (n_1722), .A (n_1345), .B (n_1344));
XOR2_X1 i_2763 (.Z (n_1721), .A (n_1396), .B (n_1395));
NOR2_X1 i_2762 (.ZN (n_1720), .A1 (n_1722), .A2 (n_1721));
AOI21_X1 i_2761 (.ZN (n_1719), .A (n_1720), .B1 (n_1722), .B2 (n_1721));
XNOR2_X1 i_2760 (.ZN (n_1718), .A (n_1324), .B (n_1317));
AOI21_X1 i_2759 (.ZN (n_1717), .A (n_1720), .B1 (n_1719), .B2 (n_1718));
XOR2_X1 i_2758 (.Z (n_1716), .A (n_1421), .B (n_1420));
XOR2_X1 i_2757 (.Z (n_1711), .A (n_1717), .B (n_1716));
XOR2_X1 i_2756 (.Z (n_1710), .A (n_1535), .B (n_1488));
XOR2_X1 i_2755 (.Z (n_1709), .A (n_1462), .B (n_1447));
XOR2_X1 i_2754 (.Z (n_1708), .A (n_1710), .B (n_1709));
XNOR2_X1 i_2753 (.ZN (n_1707), .A (n_1433), .B (n_1427));
XOR2_X1 i_2752 (.Z (n_1706), .A (n_1473), .B (n_1472));
XNOR2_X1 i_2751 (.ZN (n_1705), .A (n_1467), .B (n_1466));
XOR2_X1 i_2750 (.Z (n_1704), .A (n_1706), .B (n_1705));
XOR2_X1 i_2749 (.Z (n_1703), .A (n_1452), .B (n_1451));
NAND2_X1 i_2748 (.ZN (n_1702), .A1 (inputA[6]), .A2 (inputB[24]));
XOR2_X1 i_2747 (.Z (n_1701), .A (n_1538), .B (n_1702));
XOR2_X1 i_2746 (.Z (n_1700), .A (n_1544), .B (n_1543));
NOR2_X1 i_2745 (.ZN (n_1699), .A1 (n_1701), .A2 (n_1700));
AOI21_X1 i_2744 (.ZN (n_1698), .A (n_1699), .B1 (n_1701), .B2 (n_1700));
XNOR2_X1 i_2743 (.ZN (n_1697), .A (n_1511), .B (n_1489));
AOI22_X1 i_2742 (.ZN (n_1694), .A1 (n_1706), .A2 (n_1705), .B1 (n_1704), .B2 (n_1703));
AOI21_X1 i_2741 (.ZN (n_1693), .A (n_1699), .B1 (n_1698), .B2 (n_1697));
NAND2_X1 i_2740 (.ZN (n_1692), .A1 (n_1694), .A2 (n_1693));
OAI21_X1 i_2739 (.ZN (n_1689), .A (n_1692), .B1 (n_1694), .B2 (n_1693));
NAND2_X1 i_2738 (.ZN (n_1685), .A1 (inputA[24]), .A2 (inputB[6]));
XOR2_X1 i_2737 (.Z (n_1684), .A (n_1436), .B (n_1685));
NAND2_X1 i_2736 (.ZN (n_1682), .A1 (inputA[21]), .A2 (inputB[9]));
XOR2_X1 i_2735 (.Z (n_1681), .A (n_1440), .B (n_1682));
XNOR2_X1 i_2734 (.ZN (n_1680), .A (n_1684), .B (n_1681));
XOR2_X1 i_2733 (.Z (n_1679), .A (n_1429), .B (n_1428));
OAI22_X1 i_2732 (.ZN (n_1678), .A1 (n_1684), .A2 (n_1681), .B1 (n_1680), .B2 (n_1679));
AOI22_X1 i_2731 (.ZN (n_1677), .A1 (n_1710), .A2 (n_1709), .B1 (n_1708), .B2 (n_1707));
OAI21_X1 i_2730 (.ZN (n_1664), .A (n_1692), .B1 (n_1689), .B2 (n_1678));
INV_X1 i_2729 (.ZN (n_1663), .A (n_1664));
NOR2_X1 i_2728 (.ZN (n_1662), .A1 (n_1677), .A2 (n_1663));
AOI21_X1 i_2727 (.ZN (n_1661), .A (n_1662), .B1 (n_1677), .B2 (n_1663));
XNOR2_X1 i_2726 (.ZN (n_1660), .A (n_1416), .B (n_1413));
AOI21_X1 i_2725 (.ZN (n_1653), .A (n_1662), .B1 (n_1661), .B2 (n_1660));
AOI22_X1 i_2724 (.ZN (n_1652), .A1 (n_1717), .A2 (n_1716), .B1 (n_1711), .B2 (n_1653));
XOR2_X1 i_2723 (.Z (n_1651), .A (n_1419), .B (n_1391));
NOR2_X1 i_2722 (.ZN (n_1650), .A1 (n_1652), .A2 (n_1651));
AOI21_X1 i_2721 (.ZN (n_1649), .A (n_1650), .B1 (n_1652), .B2 (n_1651));
XNOR2_X1 i_2720 (.ZN (n_1648), .A (n_1442), .B (n_1425));
NAND2_X1 i_2719 (.ZN (n_1647), .A1 (inputA[5]), .A2 (inputB[23]));
NAND2_X1 i_2718 (.ZN (n_1646), .A1 (inputA[4]), .A2 (inputB[24]));
XNOR2_X1 i_2717 (.ZN (n_1645), .A (n_1647), .B (n_1646));
NAND2_X1 i_2716 (.ZN (n_1644), .A1 (inputA[3]), .A2 (inputB[25]));
NAND2_X1 i_2715 (.ZN (n_1643), .A1 (n_3391), .A2 (n_1301));
AOI21_X1 i_2714 (.ZN (n_1642), .A (n_22), .B1 (n_3391), .B2 (n_1301));
OAI21_X1 i_2713 (.ZN (n_1641), .A (n_1643), .B1 (n_22), .B2 (n_3097));
OAI22_X1 i_2712 (.ZN (n_1640), .A1 (n_1647), .A2 (n_1646), .B1 (n_1645), .B2 (n_1644));
XOR2_X1 i_2711 (.Z (n_1639), .A (n_1641), .B (n_1640));
NAND2_X1 i_2710 (.ZN (n_1638), .A1 (inputA[2]), .A2 (inputB[26]));
INV_X1 i_2709 (.ZN (n_1637), .A (n_1638));
AND2_X1 i_2708 (.ZN (n_1636), .A1 (inputA[1]), .A2 (inputB[27]));
NAND2_X1 i_2707 (.ZN (n_1635), .A1 (n_1637), .A2 (n_1636));
OAI21_X1 i_2706 (.ZN (n_1634), .A (n_1635), .B1 (n_1637), .B2 (n_1636));
NAND2_X1 i_2705 (.ZN (n_1633), .A1 (inputA[0]), .A2 (inputB[28]));
OAI21_X1 i_2704 (.ZN (n_1607), .A (n_1635), .B1 (n_1634), .B2 (n_1633));
AOI22_X1 i_2703 (.ZN (n_1606), .A1 (n_1641), .A2 (n_1640), .B1 (n_1639), .B2 (n_1607));
NAND2_X1 i_2702 (.ZN (n_1605), .A1 (inputA[2]), .A2 (inputB[27]));
NOR2_X1 i_2701 (.ZN (n_1604), .A1 (n_1515), .A2 (n_1605));
OAI21_X1 i_2700 (.ZN (n_1603), .A (n_23), .B1 (n_24), .B2 (n_25));
INV_X1 i_2699 (.ZN (n_1600), .A (n_1603));
NOR2_X1 i_2698 (.ZN (n_1599), .A1 (n_66), .A2 (n_128));
NOR2_X1 i_2697 (.ZN (n_1598), .A1 (n_1543), .A2 (n_1646));
AOI22_X1 i_2696 (.ZN (n_1597), .A1 (inputA[4]), .A2 (inputB[25]), .B1 (inputA[5]), .B2 (inputB[24]));
NOR2_X1 i_2695 (.ZN (n_1595), .A1 (n_1598), .A2 (n_1597));
AND2_X1 i_2694 (.ZN (n_1594), .A1 (inputA[3]), .A2 (inputB[26]));
AOI21_X1 i_2693 (.ZN (n_1593), .A (n_1604), .B1 (n_1600), .B2 (n_1599));
AOI21_X1 i_2692 (.ZN (n_1592), .A (n_1598), .B1 (n_1595), .B2 (n_1594));
XNOR2_X1 i_2691 (.ZN (n_1591), .A (n_1593), .B (n_1592));
OAI22_X1 i_2690 (.ZN (n_1586), .A1 (n_1593), .A2 (n_1592), .B1 (n_1606), .B2 (n_1591));
NAND2_X1 i_2689 (.ZN (n_1585), .A1 (inputA[5]), .A2 (inputB[27]));
NOR2_X1 i_2688 (.ZN (n_1582), .A1 (n_1546), .A2 (n_1585));
AOI22_X1 i_2687 (.ZN (n_1581), .A1 (inputA[5]), .A2 (inputB[26]), .B1 (inputA[4]), .B2 (inputB[27]));
NOR2_X1 i_2686 (.ZN (n_1580), .A1 (n_1582), .A2 (n_1581));
NAND2_X1 i_2685 (.ZN (n_1579), .A1 (inputA[0]), .A2 (inputB[31]));
XNOR2_X1 i_2684 (.ZN (n_1577), .A (n_1514), .B (n_1579));
NOR2_X1 i_2683 (.ZN (n_1576), .A1 (n_1547), .A2 (n_882));
XNOR2_X1 i_2682 (.ZN (n_1575), .A (n_833), .B (n_1580));
XOR2_X1 i_2681 (.Z (n_1574), .A (n_1577), .B (n_1576));
XOR2_X1 i_2680 (.Z (n_1573), .A (n_1575), .B (n_1574));
XOR2_X1 i_2679 (.Z (n_1572), .A (n_1211), .B (n_1210));
XOR2_X1 i_2678 (.Z (n_1571), .A (n_1185), .B (n_1184));
NAND2_X1 i_2677 (.ZN (n_1570), .A1 (n_1572), .A2 (n_1571));
OAI21_X1 i_2676 (.ZN (n_1569), .A (n_1570), .B1 (n_1572), .B2 (n_1571));
XNOR2_X1 i_2675 (.ZN (n_1568), .A (n_1332), .B (n_1327));
AOI22_X1 i_2674 (.ZN (n_1567), .A1 (n_1575), .A2 (n_1574), .B1 (n_1586), .B2 (n_1573));
OAI21_X1 i_2673 (.ZN (n_1566), .A (n_1570), .B1 (n_1569), .B2 (n_1568));
INV_X1 i_2672 (.ZN (n_1565), .A (n_1566));
NOR2_X1 i_2671 (.ZN (n_1564), .A1 (n_1567), .A2 (n_1565));
AOI21_X1 i_2670 (.ZN (n_1563), .A (n_1564), .B1 (n_1567), .B2 (n_1565));
AOI21_X1 i_2669 (.ZN (n_1562), .A (n_1564), .B1 (n_1648), .B2 (n_1563));
XNOR2_X1 i_2668 (.ZN (n_1561), .A (n_1316), .B (n_1341));
NOR2_X1 i_2667 (.ZN (n_1560), .A1 (n_1562), .A2 (n_1561));
AOI21_X1 i_2666 (.ZN (n_1559), .A (n_1560), .B1 (n_1562), .B2 (n_1561));
XNOR2_X1 i_2665 (.ZN (n_1554), .A (n_1409), .B (n_1394));
AOI21_X1 i_2664 (.ZN (n_1553), .A (n_1560), .B1 (n_1559), .B2 (n_1554));
AOI21_X1 i_2663 (.ZN (n_1552), .A (n_1650), .B1 (n_1649), .B2 (n_1553));
INV_X1 i_2662 (.ZN (n_1551), .A (inputA[8]));
INV_X1 i_2660 (.ZN (n_1547), .A (inputA[1]));
NAND2_X1 i_2659 (.ZN (n_1546), .A1 (inputA[4]), .A2 (inputB[26]));
NAND2_X1 i_2658 (.ZN (n_1545), .A1 (inputA[3]), .A2 (inputB[27]));
XNOR2_X1 i_2657 (.ZN (n_1544), .A (n_1546), .B (n_1545));
NAND2_X1 i_2656 (.ZN (n_1543), .A1 (inputA[5]), .A2 (inputB[25]));
NAND2_X1 i_2655 (.ZN (n_1542), .A1 (inputA[7]), .A2 (inputB[23]));
NAND2_X1 i_2654 (.ZN (n_1540), .A1 (inputA[8]), .A2 (inputB[22]));
XNOR2_X1 i_2653 (.ZN (n_1538), .A (n_1542), .B (n_1540));
OAI33_X1 i_2652 (.ZN (n_1537), .A1 (n_1349), .A2 (n_461), .A3 (n_1538), .B1 (n_1551)
    , .B2 (n_217), .B3 (n_1542));
OAI22_X1 i_2651 (.ZN (n_1536), .A1 (n_1546), .A2 (n_1545), .B1 (n_1544), .B2 (n_1543));
XOR2_X1 i_2650 (.Z (n_1535), .A (n_1537), .B (n_1536));
NAND2_X1 i_2649 (.ZN (n_1515), .A1 (inputA[1]), .A2 (inputB[28]));
NAND2_X1 i_2648 (.ZN (n_1514), .A1 (inputA[2]), .A2 (inputB[29]));
AOI22_X1 i_2647 (.ZN (n_1513), .A1 (inputA[1]), .A2 (inputB[29]), .B1 (inputA[2]), .B2 (inputB[28]));
INV_X1 i_2646 (.ZN (n_1512), .A (n_1513));
OAI21_X1 i_2645 (.ZN (n_1511), .A (n_1512), .B1 (n_1515), .B2 (n_1514));
NAND2_X1 i_2644 (.ZN (n_1489), .A1 (inputA[0]), .A2 (inputB[30]));
OAI22_X1 i_2643 (.ZN (n_1488), .A1 (n_1515), .A2 (n_1514), .B1 (n_1511), .B2 (n_1489));
NOR2_X1 i_2642 (.ZN (n_1487), .A1 (n_667), .A2 (n_881));
NAND3_X1 i_2641 (.ZN (n_1482), .A1 (inputA[13]), .A2 (n_1487), .A3 (inputB[18]));
INV_X1 i_2640 (.ZN (n_1480), .A (n_1482));
AOI22_X1 i_2639 (.ZN (n_1474), .A1 (inputA[13]), .A2 (inputB[17]), .B1 (inputA[12]), .B2 (inputB[18]));
NOR2_X1 i_2638 (.ZN (n_1473), .A1 (n_1480), .A2 (n_1474));
NAND2_X1 i_2637 (.ZN (n_1472), .A1 (inputA[14]), .A2 (inputB[16]));
NAND2_X1 i_2636 (.ZN (n_1471), .A1 (inputA[16]), .A2 (inputB[14]));
NAND2_X1 i_2635 (.ZN (n_1470), .A1 (inputA[17]), .A2 (inputB[13]));
XNOR2_X1 i_2634 (.ZN (n_1467), .A (n_1471), .B (n_1470));
NAND2_X1 i_2633 (.ZN (n_1466), .A1 (inputA[15]), .A2 (inputB[15]));
OAI21_X1 i_2632 (.ZN (n_1465), .A (n_1482), .B1 (n_1474), .B2 (n_1472));
OAI22_X1 i_2631 (.ZN (n_1464), .A1 (n_1471), .A2 (n_1470), .B1 (n_1467), .B2 (n_1466));
NAND2_X1 i_2630 (.ZN (n_1463), .A1 (n_1465), .A2 (n_1464));
OAI21_X1 i_2629 (.ZN (n_1462), .A (n_1463), .B1 (n_1465), .B2 (n_1464));
NAND3_X1 i_2628 (.ZN (n_1460), .A1 (inputA[10]), .A2 (n_908), .A3 (inputB[19]));
INV_X1 i_2627 (.ZN (n_1456), .A (n_1460));
AOI22_X1 i_2626 (.ZN (n_1453), .A1 (inputA[10]), .A2 (inputB[20]), .B1 (inputA[11]), .B2 (inputB[19]));
NOR2_X1 i_2625 (.ZN (n_1452), .A1 (n_1456), .A2 (n_1453));
NAND2_X1 i_2624 (.ZN (n_1451), .A1 (inputA[9]), .A2 (inputB[21]));
INV_X1 i_2623 (.ZN (n_1450), .A (n_1451));
AOI21_X1 i_2622 (.ZN (n_1447), .A (n_1456), .B1 (n_1452), .B2 (n_1450));
OAI21_X1 i_2621 (.ZN (n_1446), .A (n_1463), .B1 (n_1462), .B2 (n_1447));
INV_X1 i_2620 (.ZN (n_1445), .A (n_1446));
AOI22_X1 i_2619 (.ZN (n_1443), .A1 (n_1537), .A2 (n_1536), .B1 (n_1535), .B2 (n_1488));
XOR2_X1 i_2618 (.Z (n_1442), .A (n_1445), .B (n_1443));
NAND2_X1 i_2617 (.ZN (n_1441), .A1 (inputA[23]), .A2 (inputB[7]));
XNOR2_X1 i_2616 (.ZN (n_1440), .A (n_1209), .B (n_1441));
NAND2_X1 i_2615 (.ZN (n_1439), .A1 (inputA[26]), .A2 (inputB[4]));
XNOR2_X1 i_2614 (.ZN (n_1436), .A (n_1214), .B (n_1439));
OAI33_X1 i_2613 (.ZN (n_1435), .A1 (n_1127), .A2 (n_482), .A3 (n_1440), .B1 (n_1209)
    , .B2 (n_879), .B3 (n_213));
OAI33_X1 i_2612 (.ZN (n_1434), .A1 (n_878), .A2 (n_585), .A3 (n_1436), .B1 (n_1214)
    , .B2 (n_690), .B3 (n_214));
XOR2_X1 i_2611 (.Z (n_1433), .A (n_1435), .B (n_1434));
NAND2_X1 i_2610 (.ZN (n_1432), .A1 (inputA[19]), .A2 (inputB[10]));
NOR2_X1 i_2609 (.ZN (n_1431), .A1 (n_1199), .A2 (n_1432));
AOI22_X1 i_2608 (.ZN (n_1430), .A1 (inputA[19]), .A2 (inputB[11]), .B1 (inputA[20]), .B2 (inputB[10]));
NOR2_X1 i_2607 (.ZN (n_1429), .A1 (n_1431), .A2 (n_1430));
NOR2_X1 i_2606 (.ZN (n_1428), .A1 (n_880), .A2 (n_479));
AOI21_X1 i_2605 (.ZN (n_1427), .A (n_1431), .B1 (n_1429), .B2 (n_1428));
INV_X1 i_2604 (.ZN (n_1426), .A (n_1427));
AOI22_X1 i_2603 (.ZN (n_1425), .A1 (n_1435), .A2 (n_1434), .B1 (n_1433), .B2 (n_1426));
AOI22_X1 i_2602 (.ZN (n_1424), .A1 (n_1445), .A2 (n_1443), .B1 (n_1442), .B2 (n_1425));
XOR2_X1 i_2601 (.Z (n_1423), .A (n_821), .B (n_810));
NOR2_X1 i_2600 (.ZN (n_1422), .A1 (n_1424), .A2 (n_1423));
AOI21_X1 i_2599 (.ZN (n_1421), .A (n_1422), .B1 (n_1424), .B2 (n_1423));
XNOR2_X1 i_2598 (.ZN (n_1420), .A (n_842), .B (n_834));
AOI21_X1 i_2597 (.ZN (n_1419), .A (n_1422), .B1 (n_1421), .B2 (n_1420));
OAI21_X1 i_2596 (.ZN (n_1418), .A (n_829), .B1 (n_830), .B2 (n_858));
XOR2_X1 i_2595 (.Z (n_1417), .A (n_813), .B (n_812));
XOR2_X1 i_2594 (.Z (n_1416), .A (n_1418), .B (n_1417));
OAI21_X1 i_2593 (.ZN (n_1415), .A (inputB[30]), .B1 (n_1547), .B2 (n_129));
OAI21_X1 i_2592 (.ZN (n_1414), .A (n_921), .B1 (n_67), .B2 (n_1415));
INV_X1 i_2591 (.ZN (n_1413), .A (n_1414));
AOI22_X1 i_2590 (.ZN (n_1412), .A1 (n_1418), .A2 (n_1417), .B1 (n_1416), .B2 (n_1413));
XOR2_X1 i_2589 (.Z (n_1411), .A (n_793), .B (n_770));
NOR2_X1 i_2588 (.ZN (n_1410), .A1 (n_1412), .A2 (n_1411));
AOI21_X1 i_2587 (.ZN (n_1409), .A (n_1410), .B1 (n_1412), .B2 (n_1411));
NAND2_X1 i_2586 (.ZN (n_1408), .A1 (inputA[15]), .A2 (inputB[17]));
XNOR2_X1 i_2585 (.ZN (n_1400), .A (n_851), .B (n_1408));
OAI21_X1 i_2584 (.ZN (n_1399), .A (n_835), .B1 (n_837), .B2 (n_836));
NAND2_X1 i_2583 (.ZN (n_1398), .A1 (n_1400), .A2 (n_1399));
OAI21_X1 i_2582 (.ZN (n_1396), .A (n_1398), .B1 (n_1400), .B2 (n_1399));
XOR2_X1 i_2581 (.Z (n_1395), .A (n_826), .B (n_825));
OAI21_X1 i_2580 (.ZN (n_1394), .A (n_1398), .B1 (n_1396), .B2 (n_1395));
AOI21_X1 i_2579 (.ZN (n_1393), .A (n_1410), .B1 (n_1409), .B2 (n_1394));
XNOR2_X1 i_2578 (.ZN (n_1392), .A (n_806), .B (n_769));
XOR2_X1 i_2577 (.Z (n_1391), .A (n_1393), .B (n_1392));
AOI22_X1 i_2576 (.ZN (n_1361), .A1 (n_1393), .A2 (n_1392), .B1 (n_1419), .B2 (n_1391));
XOR2_X1 i_2575 (.Z (n_1360), .A (n_946), .B (n_944));
INV_X1 i_2574 (.ZN (n_1359), .A (n_1360));
XOR2_X1 i_2573 (.Z (n_1358), .A (n_954), .B (n_953));
INV_X1 i_2572 (.ZN (n_1357), .A (n_1358));
OAI22_X1 i_2571 (.ZN (n_1356), .A1 (n_1359), .A2 (n_1357), .B1 (n_1360), .B2 (n_1358));
INV_X1 i_2570 (.ZN (n_1355), .A (n_1356));
XOR2_X1 i_2569 (.Z (n_1350), .A (n_1361), .B (n_1356));
INV_X1 i_2568 (.ZN (n_1349), .A (inputA[6]));
INV_X1 i_2567 (.ZN (n_1348), .A (n_26));
XOR2_X1 i_2566 (.Z (n_1347), .A (n_846), .B (n_845));
XNOR2_X1 i_2565 (.ZN (n_1346), .A (n_784), .B (n_773));
XOR2_X1 i_2564 (.Z (n_1345), .A (n_1347), .B (n_1346));
XNOR2_X1 i_2563 (.ZN (n_1344), .A (n_802), .B (n_801));
AOI22_X1 i_2562 (.ZN (n_1343), .A1 (n_1347), .A2 (n_1346), .B1 (n_1345), .B2 (n_1344));
XOR2_X1 i_2561 (.Z (n_1342), .A (n_1165), .B (n_1157));
XOR2_X1 i_2560 (.Z (n_1341), .A (n_1343), .B (n_1342));
NAND2_X1 i_2559 (.ZN (n_1340), .A1 (inputB[1]), .A2 (inputA[29]));
NAND2_X1 i_2558 (.ZN (n_1339), .A1 (inputB[2]), .A2 (inputA[28]));
XNOR2_X1 i_2557 (.ZN (n_1334), .A (n_1340), .B (n_1339));
NAND2_X1 i_2556 (.ZN (n_1333), .A1 (inputB[3]), .A2 (inputA[27]));
OAI22_X1 i_2555 (.ZN (n_1332), .A1 (n_1340), .A2 (n_1339), .B1 (n_1334), .B2 (n_1333));
NOR2_X1 i_2554 (.ZN (n_1331), .A1 (n_63), .A2 (n_124));
NAND2_X1 i_2553 (.ZN (n_1330), .A1 (inputB[0]), .A2 (inputA[31]));
XOR2_X1 i_2552 (.Z (n_1327), .A (n_1331), .B (n_1330));
AOI22_X1 i_2551 (.ZN (n_1326), .A1 (n_1331), .A2 (n_1330), .B1 (n_1332), .B2 (n_1327));
XOR2_X1 i_2550 (.Z (n_1325), .A (n_1183), .B (n_1179));
XOR2_X1 i_2549 (.Z (n_1324), .A (n_1326), .B (n_1325));
XNOR2_X1 i_2548 (.ZN (n_1317), .A (n_797), .B (n_796));
AOI22_X1 i_2547 (.ZN (n_1316), .A1 (n_1326), .A2 (n_1325), .B1 (n_1324), .B2 (n_1317));
AOI22_X1 i_2546 (.ZN (n_1315), .A1 (n_1343), .A2 (n_1342), .B1 (n_1341), .B2 (n_1316));
XOR2_X1 i_2545 (.Z (n_1314), .A (n_936), .B (n_904));
NOR2_X1 i_2544 (.ZN (n_1313), .A1 (n_1315), .A2 (n_1314));
AOI21_X1 i_2543 (.ZN (n_1312), .A (n_1313), .B1 (n_1315), .B2 (n_1314));
AOI21_X1 i_2542 (.ZN (n_1311), .A (n_3279), .B1 (n_3277), .B2 (n_32));
AOI21_X1 i_2541 (.ZN (n_1310), .A (n_3284), .B1 (n_3281), .B2 (n_3280));
XNOR2_X1 i_2540 (.ZN (n_1309), .A (n_1311), .B (n_1310));
NAND2_X1 i_2539 (.ZN (n_1308), .A1 (inputB[0]), .A2 (inputA[30]));
NAND2_X1 i_2538 (.ZN (n_1307), .A1 (n_3250), .A2 (n_33));
OAI21_X1 i_2537 (.ZN (n_1306), .A (n_28), .B1 (n_29), .B2 (n_30));
NAND2_X1 i_2536 (.ZN (n_1305), .A1 (n_1307), .A2 (n_1306));
OAI21_X1 i_2535 (.ZN (n_1304), .A (n_1305), .B1 (n_1307), .B2 (n_1306));
NOR2_X1 i_2534 (.ZN (n_1303), .A1 (n_3097), .A2 (n_1542));
NOR2_X1 i_2533 (.ZN (n_1302), .A1 (n_31), .A2 (n_1303));
NOR2_X1 i_2532 (.ZN (n_1301), .A1 (n_1551), .A2 (n_216));
AOI21_X1 i_2530 (.ZN (n_1300), .A (n_1303), .B1 (n_1302), .B2 (n_1301));
OAI22_X1 i_2529 (.ZN (n_1298), .A1 (n_1311), .A2 (n_1310), .B1 (n_1309), .B2 (n_1308));
OAI21_X1 i_2528 (.ZN (n_1297), .A (n_1305), .B1 (n_1304), .B2 (n_1300));
NAND2_X1 i_2527 (.ZN (n_1296), .A1 (n_1298), .A2 (n_1297));
NOR2_X1 i_2526 (.ZN (n_1295), .A1 (n_1298), .A2 (n_1297));
AOI21_X1 i_2525 (.ZN (n_1294), .A (n_1295), .B1 (n_1298), .B2 (n_1297));
OAI22_X1 i_2524 (.ZN (n_1293), .A1 (n_3255), .A2 (n_3254), .B1 (n_3107), .B2 (n_1432));
INV_X1 i_2523 (.ZN (n_1292), .A (n_1293));
AOI21_X1 i_2522 (.ZN (n_1291), .A (n_3272), .B1 (n_3270), .B2 (n_3269));
NOR2_X1 i_2521 (.ZN (n_1290), .A1 (n_1292), .A2 (n_1291));
AOI21_X1 i_2520 (.ZN (n_1289), .A (n_1290), .B1 (n_1292), .B2 (n_1291));
OR2_X1 i_2519 (.ZN (n_1288), .A1 (n_26), .A2 (n_27));
NAND2_X1 i_2518 (.ZN (n_1287), .A1 (inputB[12]), .A2 (inputA[17]));
OAI21_X1 i_2517 (.ZN (n_1286), .A (n_1348), .B1 (n_1288), .B2 (n_1287));
AOI21_X1 i_2516 (.ZN (n_1285), .A (n_1290), .B1 (n_1289), .B2 (n_1286));
AOI21_X1 i_2515 (.ZN (n_1284), .A (n_1295), .B1 (n_1296), .B2 (n_1285));
XNOR2_X1 i_2514 (.ZN (n_1283), .A (n_924), .B (n_923));
XOR2_X1 i_2513 (.Z (n_1282), .A (n_1284), .B (n_1283));
XNOR2_X1 i_2512 (.ZN (n_1281), .A (n_911), .B (n_907));
AOI22_X1 i_2511 (.ZN (n_1280), .A1 (n_1284), .A2 (n_1283), .B1 (n_1282), .B2 (n_1281));
XOR2_X1 i_2510 (.Z (n_1254), .A (n_914), .B (n_841));
XOR2_X1 i_2509 (.Z (n_1253), .A (n_909), .B (n_908));
NOR2_X1 i_2508 (.ZN (n_1252), .A1 (n_1254), .A2 (n_1253));
AOI21_X1 i_2507 (.ZN (n_1251), .A (n_1252), .B1 (n_1254), .B2 (n_1253));
NOR2_X1 i_2506 (.ZN (n_1250), .A1 (n_1542), .A2 (n_816));
AOI22_X1 i_2505 (.ZN (n_1247), .A1 (inputB[23]), .A2 (inputA[8]), .B1 (inputB[24]), .B2 (inputA[7]));
NOR2_X1 i_2504 (.ZN (n_1246), .A1 (n_1250), .A2 (n_1247));
NOR2_X1 i_2503 (.ZN (n_1245), .A1 (n_1349), .A2 (n_219));
XNOR2_X1 i_2502 (.ZN (n_1244), .A (n_1246), .B (n_1245));
AOI21_X1 i_2501 (.ZN (n_1243), .A (n_1252), .B1 (n_1251), .B2 (n_1244));
XOR2_X1 i_2500 (.Z (n_1241), .A (n_1200), .B (n_1187));
XOR2_X1 i_2499 (.Z (n_1240), .A (n_1243), .B (n_1241));
XOR2_X1 i_2498 (.Z (n_1239), .A (n_1189), .B (n_1188));
XOR2_X1 i_2497 (.Z (n_1238), .A (n_1206), .B (n_1205));
NOR2_X1 i_2496 (.ZN (n_1232), .A1 (n_1239), .A2 (n_1238));
AOI21_X1 i_2495 (.ZN (n_1231), .A (n_1232), .B1 (n_1239), .B2 (n_1238));
XNOR2_X1 i_2494 (.ZN (n_1230), .A (n_917), .B (n_916));
AOI21_X1 i_2493 (.ZN (n_1229), .A (n_1232), .B1 (n_1231), .B2 (n_1230));
AOI22_X1 i_2492 (.ZN (n_1228), .A1 (n_1243), .A2 (n_1241), .B1 (n_1240), .B2 (n_1229));
XOR2_X1 i_2491 (.Z (n_1227), .A (n_918), .B (n_905));
XOR2_X1 i_2490 (.Z (n_1226), .A (n_1228), .B (n_1227));
AOI22_X1 i_2489 (.ZN (n_1225), .A1 (n_1228), .A2 (n_1227), .B1 (n_1280), .B2 (n_1226));
AOI21_X1 i_2488 (.ZN (n_1224), .A (n_1313), .B1 (n_1312), .B2 (n_1225));
XOR2_X1 i_2487 (.Z (n_1223), .A (n_886), .B (n_885));
XOR2_X1 i_2486 (.Z (n_1222), .A (n_1224), .B (n_1223));
XOR2_X1 i_2485 (.Z (n_1221), .A (n_1215), .B (n_1138));
AOI22_X1 i_2484 (.ZN (n_1220), .A1 (n_1224), .A2 (n_1223), .B1 (n_1222), .B2 (n_1221));
INV_X1 i_2483 (.ZN (n_1219), .A (inputB[2]));
XNOR2_X1 i_2482 (.ZN (n_1217), .A (n_1079), .B (n_1050));
XOR2_X1 i_2481 (.Z (n_1216), .A (n_747), .B (n_723));
XOR2_X1 i_2480 (.Z (n_1215), .A (n_1217), .B (n_1216));
NAND2_X1 i_2479 (.ZN (n_1214), .A1 (inputB[5]), .A2 (inputA[25]));
OR3_X1 i_2478 (.ZN (n_1213), .A1 (n_878), .A2 (n_1214), .A3 (n_214));
OAI22_X1 i_2477 (.ZN (n_1212), .A1 (n_878), .A2 (n_483), .B1 (n_214), .B2 (n_668));
NAND2_X1 i_2476 (.ZN (n_1211), .A1 (n_1213), .A2 (n_1212));
NAND2_X1 i_2475 (.ZN (n_1210), .A1 (inputB[7]), .A2 (inputA[24]));
NAND2_X1 i_2474 (.ZN (n_1209), .A1 (inputB[8]), .A2 (inputA[22]));
NOR2_X1 i_2473 (.ZN (n_1208), .A1 (n_792), .A2 (n_1209));
AOI22_X1 i_2472 (.ZN (n_1207), .A1 (inputB[9]), .A2 (inputA[22]), .B1 (inputB[8]), .B2 (inputA[23]));
NOR2_X1 i_2471 (.ZN (n_1206), .A1 (n_1208), .A2 (n_1207));
NOR2_X1 i_2470 (.ZN (n_1205), .A1 (n_1131), .A2 (n_482));
OAI21_X1 i_2469 (.ZN (n_1204), .A (n_1213), .B1 (n_1211), .B2 (n_1210));
INV_X1 i_2468 (.ZN (n_1203), .A (n_1204));
AOI21_X1 i_2467 (.ZN (n_1202), .A (n_1208), .B1 (n_1206), .B2 (n_1205));
NOR2_X1 i_2466 (.ZN (n_1201), .A1 (n_1203), .A2 (n_1202));
AOI21_X1 i_2465 (.ZN (n_1200), .A (n_1201), .B1 (n_1203), .B2 (n_1202));
NAND2_X1 i_2464 (.ZN (n_1199), .A1 (inputB[11]), .A2 (inputA[20]));
INV_X1 i_2463 (.ZN (n_1198), .A (n_1199));
NAND2_X1 i_2462 (.ZN (n_1190), .A1 (n_850), .A2 (n_1198));
OAI21_X1 i_2461 (.ZN (n_1189), .A (n_1190), .B1 (n_850), .B2 (n_1198));
NAND2_X1 i_2460 (.ZN (n_1188), .A1 (inputB[13]), .A2 (inputA[18]));
OAI21_X1 i_2459 (.ZN (n_1187), .A (n_1190), .B1 (n_1189), .B2 (n_1188));
NAND2_X1 i_2458 (.ZN (n_1186), .A1 (inputB[2]), .A2 (inputA[29]));
XNOR2_X1 i_2457 (.ZN (n_1185), .A (n_800), .B (n_1186));
NAND2_X1 i_2456 (.ZN (n_1184), .A1 (inputB[4]), .A2 (inputA[27]));
OAI22_X1 i_2455 (.ZN (n_1183), .A1 (n_800), .A2 (n_1186), .B1 (n_1185), .B2 (n_1184));
NOR2_X1 i_2454 (.ZN (n_1182), .A1 (n_1219), .A2 (n_124));
NAND2_X1 i_2453 (.ZN (n_1181), .A1 (inputB[1]), .A2 (inputA[31]));
NAND2_X1 i_2452 (.ZN (n_1180), .A1 (n_1182), .A2 (n_1181));
OAI21_X1 i_2451 (.ZN (n_1179), .A (n_1180), .B1 (n_1182), .B2 (n_1181));
INV_X1 i_2450 (.ZN (n_1169), .A (n_1179));
AOI21_X1 i_2449 (.ZN (n_1168), .A (n_1201), .B1 (n_1200), .B2 (n_1187));
AOI22_X1 i_2448 (.ZN (n_1167), .A1 (n_1182), .A2 (n_1181), .B1 (n_1183), .B2 (n_1169));
NOR2_X1 i_2447 (.ZN (n_1166), .A1 (n_1168), .A2 (n_1167));
AOI21_X1 i_2446 (.ZN (n_1165), .A (n_1166), .B1 (n_1168), .B2 (n_1167));
XOR2_X1 i_2445 (.Z (n_1157), .A (n_684), .B (n_686));
AOI21_X1 i_2444 (.ZN (n_1152), .A (n_1166), .B1 (n_1165), .B2 (n_1157));
INV_X1 i_2443 (.ZN (n_1151), .A (n_1152));
OAI21_X1 i_2442 (.ZN (n_1150), .A (n_1077), .B1 (n_1078), .B2 (n_1126));
XNOR2_X1 i_2441 (.ZN (n_1149), .A (n_1061), .B (n_1060));
XOR2_X1 i_2440 (.Z (n_1148), .A (n_1150), .B (n_1149));
XNOR2_X1 i_2439 (.ZN (n_1147), .A (n_1056), .B (n_1055));
NAND2_X1 i_2438 (.ZN (n_1146), .A1 (n_1148), .A2 (n_1147));
OAI21_X1 i_2437 (.ZN (n_1145), .A (n_744), .B1 (n_745), .B2 (n_638));
XNOR2_X1 i_2436 (.ZN (n_1144), .A (n_741), .B (n_805));
XOR2_X1 i_2435 (.Z (n_1143), .A (n_1145), .B (n_1144));
OAI21_X1 i_2434 (.ZN (n_1142), .A (n_727), .B1 (n_728), .B2 (n_849));
OAI21_X1 i_2433 (.ZN (n_1141), .A (n_1146), .B1 (n_1150), .B2 (n_1149));
AOI22_X1 i_2432 (.ZN (n_1140), .A1 (n_1145), .A2 (n_1144), .B1 (n_1143), .B2 (n_1142));
XOR2_X1 i_2431 (.Z (n_1139), .A (n_1141), .B (n_1140));
AOI22_X1 i_2430 (.ZN (n_1138), .A1 (n_1141), .A2 (n_1140), .B1 (n_1151), .B2 (n_1139));
AOI22_X1 i_2429 (.ZN (n_1137), .A1 (n_1217), .A2 (n_1216), .B1 (n_1215), .B2 (n_1138));
INV_X1 i_2428 (.ZN (n_1136), .A (inputA[11]));
INV_X1 i_2427 (.ZN (n_1132), .A (inputA[4]));
INV_X1 i_2426 (.ZN (n_1131), .A (inputB[10]));
INV_X1 i_2425 (.ZN (n_1127), .A (inputB[9]));
INV_X1 i_2424 (.ZN (n_1126), .A (n_655));
INV_X1 i_2423 (.ZN (n_1124), .A (n_767));
INV_X1 i_2422 (.ZN (n_1123), .A (n_34));
OR2_X1 i_2421 (.ZN (n_1122), .A1 (n_859), .A2 (n_128));
AND2_X1 i_2420 (.ZN (n_1112), .A1 (inputA[3]), .A2 (inputB[31]));
OR2_X1 i_2419 (.ZN (n_1109), .A1 (n_1132), .A2 (n_882));
XNOR2_X1 i_2418 (.ZN (n_1103), .A (n_1122), .B (n_1112));
OAI22_X1 i_2417 (.ZN (n_1102), .A1 (n_1122), .A2 (n_1112), .B1 (n_1109), .B2 (n_1103));
NAND2_X1 i_2416 (.ZN (n_1101), .A1 (inputA[10]), .A2 (inputB[23]));
XNOR2_X1 i_2415 (.ZN (n_1100), .A (n_631), .B (n_1101));
NAND2_X1 i_2414 (.ZN (n_1099), .A1 (inputA[8]), .A2 (inputB[25]));
OAI22_X1 i_2413 (.ZN (n_1098), .A1 (n_631), .A2 (n_1101), .B1 (n_1100), .B2 (n_1099));
INV_X1 i_2412 (.ZN (n_1097), .A (n_1098));
NAND2_X1 i_2411 (.ZN (n_1096), .A1 (inputA[6]), .A2 (inputB[27]));
XNOR2_X1 i_2410 (.ZN (n_1095), .A (n_599), .B (n_1096));
OAI33_X1 i_2409 (.ZN (n_1094), .A1 (n_859), .A2 (n_127), .A3 (n_1095), .B1 (n_812)
    , .B2 (n_864), .B3 (n_126));
INV_X1 i_2408 (.ZN (n_1093), .A (n_1094));
NAND2_X1 i_2407 (.ZN (n_1086), .A1 (inputA[3]), .A2 (inputB[30]));
XNOR2_X1 i_2406 (.ZN (n_1085), .A (n_832), .B (n_1086));
NOR2_X1 i_2405 (.ZN (n_1084), .A1 (n_67), .A2 (n_129));
OAI22_X1 i_2404 (.ZN (n_1083), .A1 (n_832), .A2 (n_1086), .B1 (n_1085), .B2 (n_1084));
INV_X1 i_2403 (.ZN (n_1082), .A (n_1083));
OAI22_X1 i_2402 (.ZN (n_1081), .A1 (n_1097), .A2 (n_1093), .B1 (n_1098), .B2 (n_1094));
OAI22_X1 i_2401 (.ZN (n_1080), .A1 (n_1097), .A2 (n_1093), .B1 (n_1082), .B2 (n_1081));
XOR2_X1 i_2400 (.Z (n_1079), .A (n_1102), .B (n_1080));
AOI21_X1 i_2399 (.ZN (n_1078), .A (n_47), .B1 (n_836), .B2 (n_650));
NAND2_X1 i_2398 (.ZN (n_1077), .A1 (n_1126), .A2 (n_1078));
NOR3_X1 i_2397 (.ZN (n_1076), .A1 (n_845), .A2 (n_480), .A3 (n_587));
AOI22_X1 i_2396 (.ZN (n_1075), .A1 (inputA[19]), .A2 (inputB[14]), .B1 (inputA[18]), .B2 (inputB[15]));
NOR2_X1 i_2395 (.ZN (n_1061), .A1 (n_1076), .A2 (n_1075));
AND2_X1 i_2394 (.ZN (n_1060), .A1 (inputA[17]), .A2 (inputB[16]));
NAND2_X1 i_2393 (.ZN (n_1059), .A1 (inputA[12]), .A2 (inputB[21]));
NOR2_X1 i_2392 (.ZN (n_1058), .A1 (n_607), .A2 (n_1059));
AOI21_X1 i_2391 (.ZN (n_1057), .A (n_1058), .B1 (n_607), .B2 (n_1059));
INV_X1 i_2390 (.ZN (n_1056), .A (n_1057));
NOR2_X1 i_2389 (.ZN (n_1055), .A1 (n_1136), .A2 (n_217));
AOI22_X1 i_2388 (.ZN (n_1054), .A1 (n_836), .A2 (n_650), .B1 (n_1126), .B2 (n_1078));
AOI21_X1 i_2387 (.ZN (n_1053), .A (n_1076), .B1 (n_1061), .B2 (n_1060));
XNOR2_X1 i_2386 (.ZN (n_1052), .A (n_1054), .B (n_1053));
AOI21_X1 i_2385 (.ZN (n_1051), .A (n_1058), .B1 (n_1057), .B2 (n_1055));
OAI22_X1 i_2384 (.ZN (n_1050), .A1 (n_1054), .A2 (n_1053), .B1 (n_1052), .B2 (n_1051));
AOI22_X1 i_2383 (.ZN (n_1049), .A1 (n_1102), .A2 (n_1080), .B1 (n_1079), .B2 (n_1050));
OAI22_X1 i_2382 (.ZN (n_1048), .A1 (n_762), .A2 (n_761), .B1 (n_598), .B2 (n_763));
NAND2_X1 i_2381 (.ZN (n_1047), .A1 (inputA[12]), .A2 (inputB[24]));
AOI22_X1 i_2380 (.ZN (n_1046), .A1 (inputA[11]), .A2 (inputB[24]), .B1 (inputA[12]), .B2 (inputB[23]));
INV_X1 i_2379 (.ZN (n_1045), .A (n_1046));
OAI21_X1 i_2378 (.ZN (n_1044), .A (n_1045), .B1 (n_610), .B2 (n_1047));
OAI22_X1 i_2377 (.ZN (n_1043), .A1 (n_610), .A2 (n_1047), .B1 (n_630), .B2 (n_1044));
XOR2_X1 i_2375 (.Z (n_1041), .A (n_1048), .B (n_1043));
AOI22_X1 i_2374 (.ZN (n_1040), .A1 (n_1124), .A2 (n_766), .B1 (n_765), .B2 (n_764));
XNOR2_X1 i_2373 (.ZN (n_1039), .A (n_1041), .B (n_1040));
XNOR2_X1 i_2372 (.ZN (n_1038), .A (n_1049), .B (n_1039));
OR2_X1 i_2371 (.ZN (n_1037), .A1 (n_217), .A2 (n_529));
XNOR2_X1 i_2370 (.ZN (n_1036), .A (n_606), .B (n_1037));
NAND2_X1 i_2369 (.ZN (n_1035), .A1 (inputA[15]), .A2 (inputB[20]));
OAI22_X1 i_2368 (.ZN (n_1029), .A1 (n_606), .A2 (n_1037), .B1 (n_1036), .B2 (n_1035));
NAND2_X1 i_2367 (.ZN (n_1028), .A1 (inputA[21]), .A2 (inputB[15]));
AOI22_X1 i_2366 (.ZN (n_1027), .A1 (inputA[20]), .A2 (inputB[15]), .B1 (inputA[21]), .B2 (inputB[14]));
INV_X1 i_2365 (.ZN (n_1026), .A (n_1027));
OAI21_X1 i_2364 (.ZN (n_1025), .A (n_1026), .B1 (n_662), .B2 (n_1028));
OAI22_X1 i_2363 (.ZN (n_1024), .A1 (n_662), .A2 (n_1028), .B1 (n_666), .B2 (n_1025));
NAND2_X1 i_2362 (.ZN (n_1023), .A1 (inputA[18]), .A2 (inputB[17]));
XNOR2_X1 i_2361 (.ZN (n_1022), .A (n_654), .B (n_1023));
OAI33_X1 i_2360 (.ZN (n_1021), .A1 (n_865), .A2 (n_314), .A3 (n_1022), .B1 (n_654)
    , .B2 (n_881), .B3 (n_479));
XOR2_X1 i_2359 (.Z (n_1020), .A (n_1024), .B (n_1021));
XOR2_X1 i_2358 (.Z (n_1019), .A (n_1029), .B (n_1020));
XOR2_X1 i_2357 (.Z (n_1018), .A (n_1038), .B (n_1019));
INV_X1 i_2356 (.ZN (n_1017), .A (n_1018));
NAND2_X1 i_2355 (.ZN (n_1016), .A1 (inputA[23]), .A2 (inputB[13]));
NAND2_X1 i_2354 (.ZN (n_1015), .A1 (inputA[24]), .A2 (inputB[11]));
NOR2_X1 i_2353 (.ZN (n_1012), .A1 (n_660), .A2 (n_1016));
AOI22_X1 i_2352 (.ZN (n_1011), .A1 (inputA[22]), .A2 (inputB[13]), .B1 (inputA[23]), .B2 (inputB[12]));
OR2_X1 i_2351 (.ZN (n_1010), .A1 (n_1012), .A2 (n_1011));
NOR2_X1 i_2350 (.ZN (n_1009), .A1 (n_1015), .A2 (n_1010));
OR2_X1 i_2349 (.ZN (n_1008), .A1 (n_1012), .A2 (n_1009));
OAI21_X1 i_2348 (.ZN (n_1007), .A (n_755), .B1 (n_752), .B2 (n_751));
NAND2_X1 i_2347 (.ZN (n_1006), .A1 (n_1008), .A2 (n_1007));
OAI21_X1 i_2346 (.ZN (n_1005), .A (n_1006), .B1 (n_1008), .B2 (n_1007));
NOR4_X1 i_2345 (.ZN (n_1004), .A1 (n_1127), .A2 (n_669), .A3 (n_214), .A4 (n_215));
AOI22_X1 i_2344 (.ZN (n_1003), .A1 (inputA[26]), .A2 (inputB[9]), .B1 (inputA[27]), .B2 (inputB[8]));
OR2_X1 i_2343 (.ZN (n_1002), .A1 (n_1004), .A2 (n_1003));
OR2_X1 i_2342 (.ZN (n_1001), .A1 (n_1131), .A2 (n_483));
NOR2_X1 i_2341 (.ZN (n_1000), .A1 (n_1002), .A2 (n_1001));
NOR2_X1 i_2340 (.ZN (n_999), .A1 (n_1004), .A2 (n_1000));
XNOR2_X1 i_2339 (.ZN (n_998), .A (n_1005), .B (n_999));
XOR2_X1 i_2338 (.Z (n_997), .A (n_1036), .B (n_1035));
NAND2_X1 i_2337 (.ZN (n_989), .A1 (inputA[16]), .A2 (inputB[19]));
XOR2_X1 i_2336 (.Z (n_983), .A (n_1022), .B (n_989));
NOR2_X1 i_2335 (.ZN (n_957), .A1 (n_997), .A2 (n_983));
AOI21_X1 i_2334 (.ZN (n_954), .A (n_957), .B1 (n_997), .B2 (n_983));
XNOR2_X1 i_2333 (.ZN (n_953), .A (n_630), .B (n_1044));
AOI21_X1 i_2332 (.ZN (n_952), .A (n_957), .B1 (n_954), .B2 (n_953));
XOR2_X1 i_2331 (.Z (n_951), .A (n_998), .B (n_952));
AOI21_X1 i_2330 (.ZN (n_950), .A (n_1000), .B1 (n_1002), .B2 (n_1001));
AOI21_X1 i_2329 (.ZN (n_949), .A (n_1009), .B1 (n_1015), .B2 (n_1010));
NOR2_X1 i_2328 (.ZN (n_948), .A1 (n_950), .A2 (n_949));
AOI21_X1 i_2327 (.ZN (n_946), .A (n_948), .B1 (n_950), .B2 (n_949));
XNOR2_X1 i_2326 (.ZN (n_944), .A (n_666), .B (n_1025));
AOI21_X1 i_2325 (.ZN (n_943), .A (n_948), .B1 (n_946), .B2 (n_944));
XOR2_X1 i_2324 (.Z (n_942), .A (n_951), .B (n_943));
XOR2_X1 i_2323 (.Z (n_941), .A (n_1018), .B (n_942));
INV_X1 i_2322 (.ZN (n_940), .A (n_941));
XOR2_X1 i_2321 (.Z (n_939), .A (n_1082), .B (n_1081));
XOR2_X1 i_2320 (.Z (n_938), .A (n_1109), .B (n_1103));
NAND2_X1 i_2319 (.ZN (n_937), .A1 (n_939), .A2 (n_938));
OAI21_X1 i_2318 (.ZN (n_936), .A (n_937), .B1 (n_939), .B2 (n_938));
AOI21_X1 i_2317 (.ZN (n_935), .A (n_1250), .B1 (n_1246), .B2 (n_1245));
AOI21_X1 i_2316 (.ZN (n_929), .A (n_1582), .B1 (n_1580), .B2 (n_40));
NOR2_X1 i_2315 (.ZN (n_925), .A1 (n_935), .A2 (n_929));
AOI21_X1 i_2314 (.ZN (n_924), .A (n_925), .B1 (n_935), .B2 (n_929));
AOI22_X1 i_2313 (.ZN (n_923), .A1 (n_41), .A2 (n_1579), .B1 (n_1577), .B2 (n_1576));
INV_X1 i_2312 (.ZN (n_922), .A (n_923));
OAI211_X1 i_2311 (.ZN (n_921), .A (inputB[31]), .B (inputA[1]), .C1 (n_882), .C2 (n_67));
INV_X1 i_2310 (.ZN (n_920), .A (n_921));
AOI21_X1 i_2309 (.ZN (n_919), .A (n_925), .B1 (n_924), .B2 (n_922));
XOR2_X1 i_2308 (.Z (n_918), .A (n_920), .B (n_919));
OR2_X1 i_2307 (.ZN (n_917), .A1 (n_34), .A2 (n_35));
NAND2_X1 i_2306 (.ZN (n_916), .A1 (inputA[15]), .A2 (inputB[16]));
NAND3_X1 i_2304 (.ZN (n_915), .A1 (inputA[13]), .A2 (n_836), .A3 (inputB[17]));
NAND2_X1 i_2303 (.ZN (n_914), .A1 (n_37), .A2 (n_915));
OAI21_X1 i_2302 (.ZN (n_913), .A (n_1123), .B1 (n_917), .B2 (n_916));
OAI21_X1 i_2301 (.ZN (n_912), .A (n_915), .B1 (n_841), .B2 (n_914));
XOR2_X1 i_2300 (.Z (n_911), .A (n_913), .B (n_912));
NOR2_X1 i_2299 (.ZN (n_910), .A1 (n_1451), .A2 (n_828));
NOR2_X1 i_2298 (.ZN (n_909), .A1 (n_38), .A2 (n_910));
NOR2_X1 i_2297 (.ZN (n_908), .A1 (n_1136), .A2 (n_414));
AOI21_X1 i_2296 (.ZN (n_907), .A (n_910), .B1 (n_909), .B2 (n_908));
INV_X1 i_2295 (.ZN (n_906), .A (n_907));
AOI22_X1 i_2294 (.ZN (n_905), .A1 (n_913), .A2 (n_912), .B1 (n_911), .B2 (n_906));
AOI22_X1 i_2293 (.ZN (n_904), .A1 (n_920), .A2 (n_919), .B1 (n_918), .B2 (n_905));
INV_X1 i_2292 (.ZN (n_903), .A (n_904));
XOR2_X1 i_2291 (.Z (n_902), .A (n_1052), .B (n_1051));
XOR2_X1 i_2290 (.Z (n_901), .A (n_731), .B (n_726));
NAND2_X1 i_2289 (.ZN (n_900), .A1 (n_902), .A2 (n_901));
OAI21_X1 i_2288 (.ZN (n_899), .A (n_900), .B1 (n_902), .B2 (n_901));
XOR2_X1 i_2287 (.Z (n_898), .A (n_1085), .B (n_1084));
XOR2_X1 i_2286 (.Z (n_897), .A (n_1100), .B (n_1099));
NOR2_X1 i_2285 (.ZN (n_896), .A1 (n_898), .A2 (n_897));
AOI21_X1 i_2284 (.ZN (n_895), .A (n_896), .B1 (n_898), .B2 (n_897));
NAND2_X1 i_2283 (.ZN (n_894), .A1 (inputA[5]), .A2 (inputB[28]));
XNOR2_X1 i_2282 (.ZN (n_893), .A (n_1095), .B (n_894));
AOI21_X1 i_2281 (.ZN (n_892), .A (n_896), .B1 (n_895), .B2 (n_893));
INV_X1 i_2280 (.ZN (n_891), .A (n_892));
OAI21_X1 i_2279 (.ZN (n_890), .A (n_937), .B1 (n_936), .B2 (n_903));
OAI21_X1 i_2278 (.ZN (n_889), .A (n_900), .B1 (n_899), .B2 (n_891));
NAND2_X1 i_2277 (.ZN (n_888), .A1 (n_890), .A2 (n_889));
INV_X1 i_2276 (.ZN (n_887), .A (n_888));
OAI21_X1 i_2275 (.ZN (n_886), .A (n_888), .B1 (n_890), .B2 (n_889));
XOR2_X1 i_2274 (.Z (n_885), .A (n_768), .B (n_758));
OAI22_X1 i_2273 (.ZN (n_884), .A1 (n_890), .A2 (n_889), .B1 (n_887), .B2 (n_885));
XOR2_X1 i_2272 (.Z (n_883), .A (n_941), .B (n_884));
INV_X1 i_2271 (.ZN (n_882), .A (inputB[30]));
INV_X1 i_2270 (.ZN (n_881), .A (inputB[17]));
INV_X1 i_2269 (.ZN (n_880), .A (inputB[12]));
INV_X1 i_2268 (.ZN (n_879), .A (inputB[7]));
INV_X1 i_2267 (.ZN (n_878), .A (inputB[6]));
INV_X1 i_2266 (.ZN (n_865), .A (inputA[16]));
INV_X1 i_2265 (.ZN (n_864), .A (inputA[7]));
INV_X1 i_2264 (.ZN (n_859), .A (inputA[5]));
INV_X1 i_2263 (.ZN (n_858), .A (n_1585));
INV_X1 i_2262 (.ZN (n_857), .A (n_688));
INV_X1 i_2260 (.ZN (n_855), .A (n_649));
INV_X1 i_2259 (.ZN (n_854), .A (n_632));
NAND2_X1 i_2258 (.ZN (n_853), .A1 (inputB[15]), .A2 (inputA[17]));
NAND2_X1 i_2257 (.ZN (n_852), .A1 (inputB[16]), .A2 (inputA[16]));
XNOR2_X1 i_2256 (.ZN (n_851), .A (n_853), .B (n_852));
NOR2_X1 i_2255 (.ZN (n_850), .A1 (n_880), .A2 (n_480));
NOR2_X1 i_2254 (.ZN (n_849), .A1 (n_671), .A2 (n_481));
NAND2_X1 i_2253 (.ZN (n_848), .A1 (n_850), .A2 (n_849));
AOI22_X1 i_2252 (.ZN (n_847), .A1 (inputB[13]), .A2 (inputA[19]), .B1 (inputB[12]), .B2 (inputA[20]));
AOI21_X1 i_2251 (.ZN (n_846), .A (n_847), .B1 (n_850), .B2 (n_849));
NAND2_X1 i_2250 (.ZN (n_845), .A1 (inputB[14]), .A2 (inputA[18]));
OAI33_X1 i_2249 (.ZN (n_844), .A1 (n_881), .A2 (n_478), .A3 (n_851), .B1 (n_865), .B2 (n_588), .B3 (n_853));
OAI21_X1 i_2248 (.ZN (n_843), .A (n_848), .B1 (n_847), .B2 (n_845));
XOR2_X1 i_2247 (.Z (n_842), .A (n_844), .B (n_843));
NAND2_X1 i_2246 (.ZN (n_841), .A1 (inputB[19]), .A2 (inputA[12]));
NOR2_X1 i_2245 (.ZN (n_839), .A1 (n_607), .A2 (n_841));
AOI22_X1 i_2244 (.ZN (n_838), .A1 (inputB[20]), .A2 (inputA[12]), .B1 (inputB[19]), .B2 (inputA[13]));
NOR2_X1 i_2243 (.ZN (n_837), .A1 (n_839), .A2 (n_838));
NOR2_X1 i_2242 (.ZN (n_836), .A1 (n_530), .A2 (n_400));
NAND2_X1 i_2241 (.ZN (n_835), .A1 (n_837), .A2 (n_836));
OAI21_X1 i_2240 (.ZN (n_834), .A (n_835), .B1 (n_607), .B2 (n_841));
NAND2_X1 i_2239 (.ZN (n_833), .A1 (inputB[28]), .A2 (inputA[3]));
NAND2_X1 i_2238 (.ZN (n_832), .A1 (inputB[29]), .A2 (inputA[4]));
NOR2_X1 i_2237 (.ZN (n_831), .A1 (n_833), .A2 (n_832));
NOR2_X1 i_2236 (.ZN (n_830), .A1 (n_39), .A2 (n_831));
NAND2_X1 i_2235 (.ZN (n_829), .A1 (n_858), .A2 (n_830));
NAND2_X1 i_2234 (.ZN (n_828), .A1 (inputB[22]), .A2 (inputA[10]));
NAND2_X1 i_2233 (.ZN (n_827), .A1 (inputB[21]), .A2 (inputA[11]));
XNOR2_X1 i_2232 (.ZN (n_826), .A (n_828), .B (n_827));
NAND2_X1 i_2231 (.ZN (n_825), .A1 (inputB[23]), .A2 (inputA[9]));
OAI21_X1 i_2230 (.ZN (n_824), .A (n_829), .B1 (n_833), .B2 (n_832));
OAI22_X1 i_2229 (.ZN (n_823), .A1 (n_828), .A2 (n_827), .B1 (n_826), .B2 (n_825));
NAND2_X1 i_2228 (.ZN (n_822), .A1 (n_824), .A2 (n_823));
OAI21_X1 i_2227 (.ZN (n_821), .A (n_822), .B1 (n_824), .B2 (n_823));
NAND2_X1 i_2226 (.ZN (n_816), .A1 (inputB[24]), .A2 (inputA[8]));
INV_X1 i_2225 (.ZN (n_815), .A (n_816));
NOR2_X1 i_2224 (.ZN (n_814), .A1 (n_864), .A2 (n_219));
XOR2_X1 i_2223 (.Z (n_813), .A (n_815), .B (n_814));
NAND2_X1 i_2222 (.ZN (n_812), .A1 (inputB[26]), .A2 (inputA[6]));
INV_X1 i_2221 (.ZN (n_811), .A (n_812));
AOI22_X1 i_2220 (.ZN (n_810), .A1 (n_815), .A2 (n_814), .B1 (n_813), .B2 (n_811));
AOI22_X1 i_2219 (.ZN (n_809), .A1 (n_844), .A2 (n_843), .B1 (n_842), .B2 (n_834));
OAI21_X1 i_2218 (.ZN (n_808), .A (n_822), .B1 (n_821), .B2 (n_810));
INV_X1 i_2217 (.ZN (n_807), .A (n_808));
XOR2_X1 i_2216 (.Z (n_806), .A (n_809), .B (n_807));
NOR2_X1 i_2215 (.ZN (n_805), .A1 (n_879), .A2 (n_214));
NAND3_X1 i_2214 (.ZN (n_804), .A1 (inputB[6]), .A2 (n_805), .A3 (inputA[25]));
OAI22_X1 i_2213 (.ZN (n_803), .A1 (n_878), .A2 (n_214), .B1 (n_879), .B2 (n_483));
NAND2_X1 i_2212 (.ZN (n_802), .A1 (n_804), .A2 (n_803));
NAND2_X1 i_2211 (.ZN (n_801), .A1 (inputB[8]), .A2 (inputA[24]));
NAND2_X1 i_2210 (.ZN (n_800), .A1 (inputB[3]), .A2 (inputA[28]));
AOI22_X1 i_2209 (.ZN (n_799), .A1 (inputB[4]), .A2 (inputA[28]), .B1 (inputB[3]), .B2 (inputA[29]));
INV_X1 i_2208 (.ZN (n_798), .A (n_799));
OAI21_X1 i_2207 (.ZN (n_797), .A (n_798), .B1 (n_682), .B2 (n_800));
NAND2_X1 i_2206 (.ZN (n_796), .A1 (inputB[5]), .A2 (inputA[27]));
OAI21_X1 i_2205 (.ZN (n_795), .A (n_804), .B1 (n_802), .B2 (n_801));
OAI22_X1 i_2204 (.ZN (n_794), .A1 (n_682), .A2 (n_800), .B1 (n_797), .B2 (n_796));
XOR2_X1 i_2203 (.Z (n_793), .A (n_795), .B (n_794));
NAND2_X1 i_2202 (.ZN (n_792), .A1 (inputB[9]), .A2 (inputA[23]));
INV_X1 i_2201 (.ZN (n_787), .A (n_792));
AND2_X1 i_2200 (.ZN (n_786), .A1 (inputB[10]), .A2 (inputA[22]));
NAND2_X1 i_2199 (.ZN (n_785), .A1 (n_787), .A2 (n_786));
OAI21_X1 i_2198 (.ZN (n_784), .A (n_785), .B1 (n_787), .B2 (n_786));
NAND2_X1 i_2197 (.ZN (n_773), .A1 (inputB[11]), .A2 (inputA[21]));
OAI21_X1 i_2196 (.ZN (n_770), .A (n_785), .B1 (n_784), .B2 (n_773));
AOI22_X1 i_2195 (.ZN (n_769), .A1 (n_795), .A2 (n_794), .B1 (n_793), .B2 (n_770));
AOI22_X1 i_2194 (.ZN (n_768), .A1 (n_809), .A2 (n_807), .B1 (n_806), .B2 (n_769));
NAND2_X1 i_2193 (.ZN (n_767), .A1 (inputB[29]), .A2 (inputA[6]));
NAND2_X1 i_2192 (.ZN (n_766), .A1 (inputB[31]), .A2 (inputA[4]));
XNOR2_X1 i_2191 (.ZN (n_765), .A (n_767), .B (n_766));
NOR2_X1 i_2190 (.ZN (n_764), .A1 (n_882), .A2 (n_859));
NAND2_X1 i_2189 (.ZN (n_763), .A1 (inputB[26]), .A2 (inputA[9]));
XNOR2_X1 i_2188 (.ZN (n_762), .A (n_598), .B (n_763));
NAND2_X1 i_2187 (.ZN (n_761), .A1 (inputB[28]), .A2 (inputA[7]));
XOR2_X1 i_2186 (.Z (n_760), .A (n_765), .B (n_764));
XOR2_X1 i_2185 (.Z (n_759), .A (n_762), .B (n_761));
XOR2_X1 i_2184 (.Z (n_758), .A (n_760), .B (n_759));
AOI22_X1 i_2183 (.ZN (n_757), .A1 (n_760), .A2 (n_759), .B1 (n_768), .B2 (n_758));
NOR2_X1 i_2182 (.ZN (n_756), .A1 (n_878), .A2 (n_124));
NAND2_X1 i_2181 (.ZN (n_755), .A1 (n_645), .A2 (n_756));
AOI22_X1 i_2180 (.ZN (n_754), .A1 (inputB[6]), .A2 (inputA[29]), .B1 (inputB[5]), .B2 (inputA[30]));
INV_X1 i_2179 (.ZN (n_753), .A (n_754));
NAND2_X1 i_2178 (.ZN (n_752), .A1 (n_755), .A2 (n_753));
NAND2_X1 i_2177 (.ZN (n_751), .A1 (inputB[7]), .A2 (inputA[28]));
AOI22_X1 i_2176 (.ZN (n_750), .A1 (n_698), .A2 (n_697), .B1 (n_857), .B2 (n_689));
XNOR2_X1 i_2175 (.ZN (n_749), .A (n_752), .B (n_751));
NOR2_X1 i_2174 (.ZN (n_748), .A1 (n_750), .A2 (n_749));
AOI21_X1 i_2173 (.ZN (n_747), .A (n_748), .B1 (n_750), .B2 (n_749));
AOI22_X1 i_2172 (.ZN (n_746), .A1 (inputB[10]), .A2 (inputA[23]), .B1 (inputB[9]), .B2 (inputA[24]));
AOI21_X1 i_2171 (.ZN (n_745), .A (n_746), .B1 (n_633), .B2 (n_787));
NAND2_X1 i_2170 (.ZN (n_744), .A1 (n_638), .A2 (n_745));
NOR2_X1 i_2169 (.ZN (n_743), .A1 (n_647), .A2 (n_796));
AOI22_X1 i_2168 (.ZN (n_742), .A1 (inputB[5]), .A2 (inputA[28]), .B1 (inputB[6]), .B2 (inputA[27]));
NOR2_X1 i_2167 (.ZN (n_741), .A1 (n_743), .A2 (n_742));
AOI22_X1 i_2166 (.ZN (n_740), .A1 (n_633), .A2 (n_787), .B1 (n_638), .B2 (n_745));
AOI21_X1 i_2165 (.ZN (n_739), .A (n_743), .B1 (n_805), .B2 (n_741));
NOR2_X1 i_2163 (.ZN (n_738), .A1 (n_740), .A2 (n_739));
AOI21_X1 i_2162 (.ZN (n_731), .A (n_738), .B1 (n_740), .B2 (n_739));
NOR2_X1 i_2161 (.ZN (n_730), .A1 (n_660), .A2 (n_773));
AOI22_X1 i_2160 (.ZN (n_729), .A1 (inputB[11]), .A2 (inputA[22]), .B1 (inputB[12]), .B2 (inputA[21]));
NOR2_X1 i_2159 (.ZN (n_728), .A1 (n_730), .A2 (n_729));
NAND2_X1 i_2158 (.ZN (n_727), .A1 (n_849), .A2 (n_728));
OAI21_X1 i_2157 (.ZN (n_726), .A (n_727), .B1 (n_660), .B2 (n_773));
AOI21_X1 i_2156 (.ZN (n_723), .A (n_738), .B1 (n_731), .B2 (n_726));
INV_X1 i_2155 (.ZN (n_722), .A (n_723));
AOI21_X1 i_2154 (.ZN (n_721), .A (n_748), .B1 (n_747), .B2 (n_722));
XOR2_X1 i_2153 (.Z (n_720), .A (n_757), .B (n_721));
AOI22_X1 i_2152 (.ZN (n_719), .A1 (n_855), .A2 (n_656), .B1 (n_657), .B2 (n_661));
AOI22_X1 i_2151 (.ZN (n_717), .A1 (n_854), .A2 (n_639), .B1 (n_641), .B2 (n_640));
NOR2_X1 i_2150 (.ZN (n_716), .A1 (n_608), .A2 (n_601));
AOI21_X1 i_2149 (.ZN (n_715), .A (n_716), .B1 (n_600), .B2 (n_593));
XOR2_X1 i_2148 (.Z (n_714), .A (n_717), .B (n_715));
XOR2_X1 i_2147 (.Z (n_712), .A (n_719), .B (n_714));
INV_X1 i_2146 (.ZN (n_711), .A (n_712));
XOR2_X1 i_2145 (.Z (n_710), .A (n_720), .B (n_712));
AOI21_X1 i_2144 (.ZN (n_709), .A (n_706), .B1 (n_708), .B2 (n_707));
INV_X1 i_2143 (.ZN (n_708), .A (n_703));
AOI21_X1 i_2142 (.ZN (n_707), .A (n_706), .B1 (n_705), .B2 (n_704));
NOR2_X1 i_2141 (.ZN (n_706), .A1 (n_704), .A2 (n_705));
AOI22_X1 i_2140 (.ZN (n_705), .A1 (n_674), .A2 (n_675), .B1 (n_672), .B2 (n_673));
AOI21_X1 i_2139 (.ZN (n_704), .A (n_679), .B1 (n_680), .B2 (n_681));
AOI22_X1 i_2138 (.ZN (n_703), .A1 (n_701), .A2 (n_702), .B1 (n_699), .B2 (n_700));
XNOR2_X1 i_2137 (.ZN (n_702), .A (n_643), .B (n_642));
XOR2_X1 i_2136 (.Z (n_701), .A (n_699), .B (n_700));
XOR2_X1 i_2135 (.Z (n_700), .A (n_635), .B (n_634));
XNOR2_X1 i_2134 (.ZN (n_699), .A (n_698), .B (n_697));
XNOR2_X1 i_2133 (.ZN (n_698), .A (n_688), .B (n_689));
NOR2_X1 i_2132 (.ZN (n_697), .A1 (n_690), .A2 (n_124));
INV_X1 i_2131 (.ZN (n_690), .A (inputB[4]));
NAND2_X1 i_2130 (.ZN (n_689), .A1 (inputB[3]), .A2 (inputA[31]));
AOI22_X1 i_2129 (.ZN (n_688), .A1 (n_684), .A2 (n_686), .B1 (n_687), .B2 (n_683));
INV_X1 i_2128 (.ZN (n_687), .A (n_682));
NOR2_X1 i_2126 (.ZN (n_686), .A1 (n_685), .A2 (n_124));
INV_X1 i_2125 (.ZN (n_685), .A (inputB[3]));
XNOR2_X1 i_2124 (.ZN (n_684), .A (n_682), .B (n_683));
NAND2_X1 i_2123 (.ZN (n_683), .A1 (inputB[2]), .A2 (inputA[31]));
NAND2_X1 i_2122 (.ZN (n_682), .A1 (inputA[29]), .A2 (inputB[4]));
XNOR2_X1 i_2121 (.ZN (n_681), .A (n_651), .B (n_650));
AOI21_X1 i_2120 (.ZN (n_680), .A (n_679), .B1 (n_677), .B2 (n_678));
NOR2_X1 i_2119 (.ZN (n_679), .A1 (n_677), .A2 (n_678));
XOR2_X1 i_2118 (.Z (n_678), .A (n_663), .B (n_662));
XOR2_X1 i_2117 (.Z (n_677), .A (n_676), .B (n_658));
NAND2_X1 i_2116 (.ZN (n_676), .A1 (inputB[13]), .A2 (inputA[21]));
XNOR2_X1 i_2115 (.ZN (n_675), .A (n_595), .B (n_594));
XOR2_X1 i_2114 (.Z (n_674), .A (n_672), .B (n_673));
XNOR2_X1 i_2113 (.ZN (n_673), .A (n_603), .B (n_602));
XOR2_X1 i_2112 (.Z (n_672), .A (n_627), .B (n_610));
INV_X1 i_2111 (.ZN (n_671), .A (inputB[13]));
INV_X1 i_2110 (.ZN (n_670), .A (inputB[11]));
INV_X1 i_2109 (.ZN (n_669), .A (inputB[8]));
INV_X1 i_2108 (.ZN (n_668), .A (inputB[5]));
INV_X1 i_2107 (.ZN (n_667), .A (inputA[12]));
NAND2_X1 i_2106 (.ZN (n_666), .A1 (inputB[16]), .A2 (inputA[19]));
OR3_X1 i_2105 (.ZN (n_665), .A1 (n_587), .A2 (n_666), .A3 (n_479));
OAI22_X1 i_2104 (.ZN (n_664), .A1 (n_587), .A2 (n_480), .B1 (n_479), .B2 (n_588));
NAND2_X1 i_2103 (.ZN (n_663), .A1 (n_665), .A2 (n_664));
NAND2_X1 i_2102 (.ZN (n_662), .A1 (inputB[14]), .A2 (inputA[20]));
OAI21_X1 i_2101 (.ZN (n_661), .A (n_665), .B1 (n_663), .B2 (n_662));
NAND2_X1 i_2100 (.ZN (n_660), .A1 (inputB[12]), .A2 (inputA[22]));
NAND2_X1 i_2099 (.ZN (n_659), .A1 (inputB[11]), .A2 (inputA[23]));
XNOR2_X1 i_2098 (.ZN (n_658), .A (n_660), .B (n_659));
OAI33_X1 i_2097 (.ZN (n_657), .A1 (n_671), .A2 (n_482), .A3 (n_658), .B1 (n_670), .B2 (n_213), .B3 (n_660));
XOR2_X1 i_2096 (.Z (n_656), .A (n_661), .B (n_657));
NAND2_X1 i_2095 (.ZN (n_655), .A1 (inputB[17]), .A2 (inputA[16]));
NAND2_X1 i_2094 (.ZN (n_654), .A1 (inputB[18]), .A2 (inputA[17]));
NOR2_X1 i_2093 (.ZN (n_653), .A1 (n_655), .A2 (n_654));
AOI22_X1 i_2092 (.ZN (n_652), .A1 (inputB[17]), .A2 (inputA[17]), .B1 (inputB[18]), .B2 (inputA[16]));
NOR2_X1 i_2091 (.ZN (n_651), .A1 (n_653), .A2 (n_652));
NOR2_X1 i_2090 (.ZN (n_650), .A1 (n_478), .A2 (n_314));
AOI21_X1 i_2089 (.ZN (n_649), .A (n_653), .B1 (n_651), .B2 (n_650));
XOR2_X1 i_2088 (.Z (n_648), .A (n_656), .B (n_649));
NAND2_X1 i_2087 (.ZN (n_647), .A1 (inputB[6]), .A2 (inputA[28]));
INV_X1 i_2086 (.ZN (n_646), .A (n_647));
NOR2_X1 i_2085 (.ZN (n_645), .A1 (n_668), .A2 (n_123));
NAND2_X1 i_2084 (.ZN (n_644), .A1 (n_646), .A2 (n_645));
OAI21_X1 i_2083 (.ZN (n_643), .A (n_644), .B1 (n_646), .B2 (n_645));
NAND2_X1 i_2082 (.ZN (n_642), .A1 (inputB[7]), .A2 (inputA[27]));
OAI21_X1 i_2081 (.ZN (n_641), .A (n_644), .B1 (n_643), .B2 (n_642));
NAND2_X1 i_2080 (.ZN (n_640), .A1 (inputB[4]), .A2 (inputA[31]));
XOR2_X1 i_2079 (.Z (n_639), .A (n_641), .B (n_640));
NOR2_X1 i_2078 (.ZN (n_638), .A1 (n_669), .A2 (n_483));
AND3_X1 i_2077 (.ZN (n_637), .A1 (inputB[9]), .A2 (n_638), .A3 (inputA[26]));
AOI22_X1 i_2076 (.ZN (n_636), .A1 (inputB[8]), .A2 (inputA[26]), .B1 (inputB[9]), .B2 (inputA[25]));
NOR2_X1 i_2075 (.ZN (n_635), .A1 (n_637), .A2 (n_636));
NAND2_X1 i_2074 (.ZN (n_634), .A1 (inputB[10]), .A2 (inputA[24]));
INV_X1 i_2073 (.ZN (n_633), .A (n_634));
AOI21_X1 i_2072 (.ZN (n_632), .A (n_637), .B1 (n_635), .B2 (n_633));
NAND2_X1 i_2071 (.ZN (n_631), .A1 (inputB[24]), .A2 (inputA[9]));
NAND2_X1 i_2070 (.ZN (n_630), .A1 (inputB[25]), .A2 (inputA[10]));
NOR2_X1 i_2069 (.ZN (n_629), .A1 (n_631), .A2 (n_630));
AOI22_X1 i_2068 (.ZN (n_628), .A1 (inputB[24]), .A2 (inputA[10]), .B1 (inputB[25]), .B2 (inputA[9]));
NOR2_X1 i_2067 (.ZN (n_627), .A1 (n_629), .A2 (n_628));
NAND2_X1 i_2066 (.ZN (n_610), .A1 (inputB[23]), .A2 (inputA[11]));
INV_X1 i_2065 (.ZN (n_609), .A (n_610));
AOI21_X1 i_2064 (.ZN (n_608), .A (n_629), .B1 (n_627), .B2 (n_609));
NAND2_X1 i_2063 (.ZN (n_607), .A1 (inputB[20]), .A2 (inputA[13]));
NAND2_X1 i_2062 (.ZN (n_606), .A1 (inputB[21]), .A2 (inputA[14]));
NOR2_X1 i_2061 (.ZN (n_605), .A1 (n_607), .A2 (n_606));
AOI22_X1 i_2060 (.ZN (n_604), .A1 (inputB[21]), .A2 (inputA[13]), .B1 (inputB[20]), .B2 (inputA[14]));
NOR2_X1 i_2059 (.ZN (n_603), .A1 (n_605), .A2 (n_604));
NOR2_X1 i_2058 (.ZN (n_602), .A1 (n_667), .A2 (n_217));
AOI21_X1 i_2057 (.ZN (n_601), .A (n_605), .B1 (n_603), .B2 (n_602));
XOR2_X1 i_2056 (.Z (n_600), .A (n_608), .B (n_601));
NAND2_X1 i_2055 (.ZN (n_599), .A1 (inputB[26]), .A2 (inputA[7]));
NAND2_X1 i_2054 (.ZN (n_598), .A1 (inputB[27]), .A2 (inputA[8]));
AOI22_X1 i_2053 (.ZN (n_597), .A1 (inputB[26]), .A2 (inputA[8]), .B1 (inputB[27]), .B2 (inputA[7]));
INV_X1 i_2052 (.ZN (n_596), .A (n_597));
OAI21_X1 i_2051 (.ZN (n_595), .A (n_596), .B1 (n_599), .B2 (n_598));
NAND2_X1 i_2050 (.ZN (n_594), .A1 (inputB[28]), .A2 (inputA[6]));
OAI22_X1 i_2049 (.ZN (n_593), .A1 (n_599), .A2 (n_598), .B1 (n_595), .B2 (n_594));
XOR2_X1 i_2048 (.Z (n_592), .A (n_639), .B (n_632));
XNOR2_X1 i_2047 (.ZN (n_591), .A (n_600), .B (n_593));
XOR2_X1 i_2046 (.Z (n_590), .A (n_592), .B (n_591));
AOI22_X1 i_2045 (.ZN (n_589), .A1 (n_592), .A2 (n_591), .B1 (n_648), .B2 (n_590));
INV_X1 i_2044 (.ZN (n_588), .A (inputB[16]));
INV_X1 i_2043 (.ZN (n_587), .A (inputB[15]));
INV_X1 i_2042 (.ZN (n_586), .A (inputB[14]));
INV_X1 i_2041 (.ZN (n_585), .A (inputA[24]));
NAND2_X1 i_2040 (.ZN (n_584), .A1 (inputB[17]), .A2 (inputA[26]));
NAND2_X1 i_2039 (.ZN (n_583), .A1 (inputB[18]), .A2 (inputA[27]));
AOI22_X1 i_2038 (.ZN (n_582), .A1 (inputB[17]), .A2 (inputA[27]), .B1 (inputB[18]), .B2 (inputA[26]));
INV_X1 i_2037 (.ZN (n_581), .A (n_582));
OAI21_X1 i_2036 (.ZN (n_579), .A (n_581), .B1 (n_584), .B2 (n_583));
NAND2_X1 i_2035 (.ZN (n_578), .A1 (inputB[19]), .A2 (inputA[25]));
NAND2_X1 i_2034 (.ZN (n_577), .A1 (inputB[15]), .A2 (inputA[29]));
NAND2_X1 i_2033 (.ZN (n_576), .A1 (inputB[14]), .A2 (inputA[30]));
XNOR2_X1 i_2032 (.ZN (n_575), .A (n_577), .B (n_576));
NOR2_X1 i_2031 (.ZN (n_574), .A1 (n_587), .A2 (n_124));
OAI33_X1 i_2030 (.ZN (n_573), .A1 (n_588), .A2 (n_122), .A3 (n_575), .B1 (n_586), .B2 (n_124), .B3 (n_577));
OAI22_X1 i_2029 (.ZN (n_572), .A1 (n_584), .A2 (n_583), .B1 (n_579), .B2 (n_578));
XOR2_X1 i_2028 (.Z (n_571), .A (n_573), .B (n_572));
NAND2_X1 i_2027 (.ZN (n_570), .A1 (inputB[21]), .A2 (inputA[24]));
OR3_X1 i_2026 (.ZN (n_569), .A1 (n_414), .A2 (n_570), .A3 (n_213));
OAI22_X1 i_2025 (.ZN (n_568), .A1 (n_585), .A2 (n_414), .B1 (n_213), .B2 (n_216));
NAND2_X1 i_2024 (.ZN (n_567), .A1 (n_569), .A2 (n_568));
NAND2_X1 i_2023 (.ZN (n_566), .A1 (inputB[22]), .A2 (inputA[22]));
OAI21_X1 i_2022 (.ZN (n_565), .A (n_569), .B1 (n_567), .B2 (n_566));
NAND2_X1 i_2021 (.ZN (n_564), .A1 (n_397), .A2 (n_399));
XOR2_X1 i_2020 (.Z (n_563), .A (n_395), .B (n_564));
AOI22_X1 i_2019 (.ZN (n_562), .A1 (n_573), .A2 (n_572), .B1 (n_571), .B2 (n_565));
NAND2_X1 i_2018 (.ZN (n_561), .A1 (n_563), .A2 (n_562));
NOR2_X1 i_2017 (.ZN (n_560), .A1 (n_563), .A2 (n_562));
INV_X1 i_2016 (.ZN (n_559), .A (n_560));
NOR2_X1 i_2014 (.ZN (n_558), .A1 (n_588), .A2 (n_123));
NAND2_X1 i_2013 (.ZN (n_557), .A1 (inputB[14]), .A2 (inputA[31]));
XOR2_X1 i_2012 (.Z (n_556), .A (n_558), .B (n_557));
AOI22_X1 i_2011 (.ZN (n_555), .A1 (n_558), .A2 (n_557), .B1 (n_574), .B2 (n_556));
NAND2_X1 i_2010 (.ZN (n_554), .A1 (inputB[15]), .A2 (inputA[31]));
XNOR2_X1 i_2009 (.ZN (n_553), .A (n_555), .B (n_554));
NOR2_X1 i_2008 (.ZN (n_552), .A1 (n_588), .A2 (n_124));
XOR2_X1 i_2007 (.Z (n_551), .A (n_553), .B (n_552));
OAI21_X1 i_2006 (.ZN (n_550), .A (n_561), .B1 (n_560), .B2 (n_551));
XOR2_X1 i_2005 (.Z (n_549), .A (n_457), .B (n_276));
XOR2_X1 i_2004 (.Z (n_548), .A (n_384), .B (n_383));
NOR2_X1 i_2001 (.ZN (n_547), .A1 (n_549), .A2 (n_548));
AOI21_X1 i_2000 (.ZN (n_546), .A (n_547), .B1 (n_549), .B2 (n_548));
NAND2_X1 i_1999 (.ZN (n_545), .A1 (inputB[28]), .A2 (inputA[18]));
XNOR2_X1 i_1998 (.ZN (n_544), .A (n_451), .B (n_545));
AOI21_X1 i_1997 (.ZN (n_543), .A (n_547), .B1 (n_546), .B2 (n_544));
XOR2_X1 i_1996 (.Z (n_534), .A (n_390), .B (n_382));
NOR2_X1 i_1995 (.ZN (n_533), .A1 (n_543), .A2 (n_534));
AOI21_X1 i_1994 (.ZN (n_532), .A (n_533), .B1 (n_543), .B2 (n_534));
AOI21_X1 i_1993 (.ZN (n_531), .A (n_533), .B1 (n_550), .B2 (n_532));
INV_X1 i_1992 (.ZN (n_530), .A (inputA[14]));
INV_X1 i_1991 (.ZN (n_529), .A (inputA[13]));
XOR2_X1 i_1990 (.Z (n_528), .A (n_448), .B (n_441));
XOR2_X1 i_1989 (.Z (n_527), .A (n_438), .B (n_437));
XOR2_X1 i_1988 (.Z (n_526), .A (n_528), .B (n_527));
NAND2_X1 i_1987 (.ZN (n_525), .A1 (inputA[18]), .A2 (inputB[26]));
AOI22_X1 i_1986 (.ZN (n_524), .A1 (inputA[18]), .A2 (inputB[27]), .B1 (inputA[19]), .B2 (inputB[26]));
INV_X1 i_1985 (.ZN (n_523), .A (n_524));
OAI21_X1 i_1984 (.ZN (n_522), .A (n_523), .B1 (n_456), .B2 (n_525));
NAND2_X1 i_1983 (.ZN (n_521), .A1 (inputA[17]), .A2 (inputB[28]));
NAND2_X1 i_1982 (.ZN (n_518), .A1 (inputA[15]), .A2 (inputB[29]));
AOI22_X1 i_1981 (.ZN (n_517), .A1 (inputA[16]), .A2 (inputB[29]), .B1 (inputA[15]), .B2 (inputB[30]));
INV_X1 i_1980 (.ZN (n_516), .A (n_517));
OAI21_X1 i_1979 (.ZN (n_515), .A (n_516), .B1 (n_444), .B2 (n_518));
NOR2_X1 i_1978 (.ZN (n_514), .A1 (n_530), .A2 (n_129));
NAND2_X1 i_1977 (.ZN (n_513), .A1 (inputA[17]), .A2 (inputB[27]));
XNOR2_X1 i_1976 (.ZN (n_512), .A (n_525), .B (n_513));
NAND2_X1 i_1975 (.ZN (n_511), .A1 (inputA[16]), .A2 (inputB[28]));
NAND2_X1 i_1974 (.ZN (n_510), .A1 (inputA[19]), .A2 (inputB[24]));
NAND2_X1 i_1973 (.ZN (n_509), .A1 (inputA[20]), .A2 (inputB[25]));
NOR2_X1 i_1972 (.ZN (n_508), .A1 (n_510), .A2 (n_509));
AOI22_X1 i_1971 (.ZN (n_507), .A1 (inputA[20]), .A2 (inputB[24]), .B1 (inputA[19]), .B2 (inputB[25]));
NOR2_X1 i_1970 (.ZN (n_506), .A1 (n_508), .A2 (n_507));
NOR2_X1 i_1969 (.ZN (n_500), .A1 (n_482), .A2 (n_218));
AOI21_X1 i_1968 (.ZN (n_499), .A (n_508), .B1 (n_506), .B2 (n_500));
OAI22_X1 i_1967 (.ZN (n_498), .A1 (n_525), .A2 (n_513), .B1 (n_512), .B2 (n_511));
INV_X1 i_1966 (.ZN (n_497), .A (n_498));
NOR2_X1 i_1965 (.ZN (n_496), .A1 (n_499), .A2 (n_497));
AOI21_X1 i_1964 (.ZN (n_495), .A (n_496), .B1 (n_499), .B2 (n_497));
NAND2_X1 i_1963 (.ZN (n_494), .A1 (inputA[14]), .A2 (inputB[30]));
XNOR2_X1 i_1962 (.ZN (n_493), .A (n_518), .B (n_494));
NOR2_X1 i_1961 (.ZN (n_492), .A1 (n_529), .A2 (n_129));
OAI22_X1 i_1960 (.ZN (n_491), .A1 (n_518), .A2 (n_494), .B1 (n_493), .B2 (n_492));
AOI21_X1 i_1959 (.ZN (n_490), .A (n_496), .B1 (n_495), .B2 (n_491));
OAI22_X1 i_1958 (.ZN (n_489), .A1 (n_456), .A2 (n_525), .B1 (n_522), .B2 (n_521));
OAI22_X1 i_1957 (.ZN (n_488), .A1 (n_444), .A2 (n_518), .B1 (n_515), .B2 (n_514));
NAND2_X1 i_1956 (.ZN (n_487), .A1 (n_489), .A2 (n_488));
OAI21_X1 i_1955 (.ZN (n_486), .A (n_487), .B1 (n_489), .B2 (n_488));
OAI21_X1 i_1954 (.ZN (n_485), .A (n_487), .B1 (n_490), .B2 (n_486));
AOI22_X1 i_1953 (.ZN (n_484), .A1 (n_528), .A2 (n_527), .B1 (n_526), .B2 (n_485));
INV_X1 i_1952 (.ZN (n_483), .A (inputA[25]));
INV_X1 i_1951 (.ZN (n_482), .A (inputA[21]));
INV_X1 i_1950 (.ZN (n_481), .A (inputA[20]));
INV_X1 i_1949 (.ZN (n_480), .A (inputA[19]));
INV_X1 i_1948 (.ZN (n_479), .A (inputA[18]));
INV_X1 i_1947 (.ZN (n_478), .A (inputA[15]));
INV_X1 i_1945 (.ZN (n_461), .A (inputB[24]));
INV_X1 i_1944 (.ZN (n_460), .A (n_372));
OR3_X1 i_1943 (.ZN (n_459), .A1 (n_482), .A2 (n_271), .A3 (n_461));
OAI22_X1 i_1942 (.ZN (n_458), .A1 (n_461), .A2 (n_259), .B1 (n_482), .B2 (n_219));
NAND2_X1 i_1941 (.ZN (n_457), .A1 (n_459), .A2 (n_458));
NAND2_X1 i_1940 (.ZN (n_456), .A1 (inputA[19]), .A2 (inputB[27]));
NAND2_X1 i_1939 (.ZN (n_452), .A1 (inputA[20]), .A2 (inputB[26]));
XNOR2_X1 i_1938 (.ZN (n_451), .A (n_456), .B (n_452));
OAI21_X1 i_1937 (.ZN (n_450), .A (n_459), .B1 (n_276), .B2 (n_457));
OAI33_X1 i_1936 (.ZN (n_449), .A1 (n_480), .A2 (n_126), .A3 (n_452), .B1 (n_479), .B2 (n_127), .B3 (n_451));
XOR2_X1 i_1935 (.Z (n_448), .A (n_450), .B (n_449));
NOR2_X1 i_1934 (.ZN (n_447), .A1 (n_478), .A2 (n_129));
NAND2_X1 i_1933 (.ZN (n_446), .A1 (inputA[17]), .A2 (inputB[29]));
XOR2_X1 i_1932 (.Z (n_445), .A (n_447), .B (n_446));
NAND2_X1 i_1931 (.ZN (n_444), .A1 (inputA[16]), .A2 (inputB[30]));
INV_X1 i_1930 (.ZN (n_443), .A (n_444));
NAND2_X1 i_1929 (.ZN (n_442), .A1 (n_445), .A2 (n_443));
OAI21_X1 i_1928 (.ZN (n_441), .A (n_442), .B1 (n_447), .B2 (n_446));
AOI22_X1 i_1927 (.ZN (n_440), .A1 (n_450), .A2 (n_449), .B1 (n_448), .B2 (n_441));
AND2_X1 i_1926 (.ZN (n_439), .A1 (inputA[16]), .A2 (inputB[31]));
XNOR2_X1 i_1925 (.ZN (n_438), .A (n_268), .B (n_439));
NAND2_X1 i_1924 (.ZN (n_437), .A1 (inputA[17]), .A2 (inputB[30]));
NOR2_X1 i_1923 (.ZN (n_436), .A1 (n_330), .A2 (n_452));
AOI22_X1 i_1922 (.ZN (n_433), .A1 (inputA[20]), .A2 (inputB[27]), .B1 (inputA[21]), .B2 (inputB[26]));
NOR2_X1 i_1921 (.ZN (n_432), .A1 (n_436), .A2 (n_433));
NOR2_X1 i_1920 (.ZN (n_431), .A1 (n_480), .A2 (n_127));
AOI21_X1 i_1919 (.ZN (n_430), .A (n_436), .B1 (n_432), .B2 (n_431));
OAI22_X1 i_1918 (.ZN (n_429), .A1 (n_268), .A2 (n_439), .B1 (n_438), .B2 (n_437));
INV_X1 i_1917 (.ZN (n_428), .A (n_429));
XNOR2_X1 i_1916 (.ZN (n_427), .A (n_430), .B (n_428));
OAI22_X1 i_1915 (.ZN (n_426), .A1 (n_430), .A2 (n_428), .B1 (n_440), .B2 (n_427));
NAND2_X1 i_1914 (.ZN (n_425), .A1 (n_460), .A2 (n_360));
OAI22_X1 i_1913 (.ZN (n_424), .A1 (n_328), .A2 (n_327), .B1 (n_330), .B2 (n_329));
XOR2_X1 i_1912 (.Z (n_423), .A (n_425), .B (n_424));
OAI33_X1 i_1911 (.ZN (n_422), .A1 (n_219), .A2 (n_340), .A3 (n_213), .B1 (n_483), .B2 (n_275), .B3 (n_218));
XOR2_X1 i_1910 (.Z (n_421), .A (n_423), .B (n_422));
NOR2_X1 i_1909 (.ZN (n_420), .A1 (n_481), .A2 (n_128));
NAND2_X1 i_1908 (.ZN (n_419), .A1 (inputA[18]), .A2 (inputB[31]));
XOR2_X1 i_1907 (.Z (n_418), .A (n_420), .B (n_419));
XNOR2_X1 i_1906 (.ZN (n_417), .A (n_267), .B (n_418));
XOR2_X1 i_1905 (.Z (n_416), .A (n_421), .B (n_417));
XOR2_X1 i_1904 (.Z (n_415), .A (n_426), .B (n_416));
INV_X1 i_1903 (.ZN (n_414), .A (inputB[20]));
INV_X1 i_1902 (.ZN (n_400), .A (inputB[18]));
OAI21_X1 i_1901 (.ZN (n_399), .A (n_285), .B1 (n_400), .B2 (n_122));
NOR3_X1 i_1900 (.ZN (n_398), .A1 (n_400), .A2 (n_285), .A3 (n_122));
INV_X1 i_1899 (.ZN (n_397), .A (n_398));
NOR2_X1 i_1898 (.ZN (n_395), .A1 (n_314), .A2 (n_215));
AND2_X1 i_1897 (.ZN (n_394), .A1 (inputB[16]), .A2 (inputA[31]));
OAI21_X1 i_1896 (.ZN (n_393), .A (n_399), .B1 (n_398), .B2 (n_395));
NOR2_X1 i_1895 (.ZN (n_392), .A1 (n_394), .A2 (n_393));
AOI21_X1 i_1894 (.ZN (n_390), .A (n_392), .B1 (n_394), .B2 (n_393));
NAND2_X1 i_1893 (.ZN (n_389), .A1 (inputB[20]), .A2 (inputA[25]));
AOI22_X1 i_1892 (.ZN (n_388), .A1 (inputB[20]), .A2 (inputA[26]), .B1 (inputB[21]), .B2 (inputA[25]));
INV_X1 i_1891 (.ZN (n_385), .A (n_388));
OAI21_X1 i_1890 (.ZN (n_384), .A (n_385), .B1 (n_301), .B2 (n_389));
NAND2_X1 i_1889 (.ZN (n_383), .A1 (inputB[22]), .A2 (inputA[24]));
OAI22_X1 i_1888 (.ZN (n_382), .A1 (n_301), .A2 (n_389), .B1 (n_384), .B2 (n_383));
AOI21_X1 i_1887 (.ZN (n_381), .A (n_392), .B1 (n_390), .B2 (n_382));
XOR2_X1 i_1886 (.Z (n_376), .A (n_311), .B (n_310));
XOR2_X1 i_1885 (.Z (n_375), .A (n_381), .B (n_376));
NAND2_X1 i_1884 (.ZN (n_373), .A1 (inputB[22]), .A2 (inputA[27]));
NOR2_X1 i_1883 (.ZN (n_372), .A1 (n_301), .A2 (n_373));
NOR2_X1 i_1882 (.ZN (n_363), .A1 (n_414), .A2 (n_122));
AOI22_X1 i_1881 (.ZN (n_362), .A1 (inputB[22]), .A2 (inputA[26]), .B1 (inputB[21]), .B2 (inputA[27]));
NOR2_X1 i_1880 (.ZN (n_361), .A1 (n_372), .A2 (n_362));
NAND2_X1 i_1879 (.ZN (n_360), .A1 (n_363), .A2 (n_361));
OAI21_X1 i_1878 (.ZN (n_359), .A (n_360), .B1 (n_363), .B2 (n_361));
NAND2_X1 i_1877 (.ZN (n_358), .A1 (inputB[23]), .A2 (inputA[25]));
XNOR2_X1 i_1876 (.ZN (n_340), .A (n_275), .B (n_358));
NAND2_X1 i_1875 (.ZN (n_339), .A1 (inputB[25]), .A2 (inputA[23]));
XOR2_X1 i_1874 (.Z (n_338), .A (n_340), .B (n_339));
XOR2_X1 i_1873 (.Z (n_334), .A (n_264), .B (n_263));
NOR2_X1 i_1872 (.ZN (n_333), .A1 (n_338), .A2 (n_334));
AOI21_X1 i_1871 (.ZN (n_331), .A (n_333), .B1 (n_338), .B2 (n_334));
NAND2_X1 i_1870 (.ZN (n_330), .A1 (inputB[27]), .A2 (inputA[21]));
NAND2_X1 i_1869 (.ZN (n_329), .A1 (inputB[26]), .A2 (inputA[22]));
XNOR2_X1 i_1868 (.ZN (n_328), .A (n_330), .B (n_329));
NAND2_X1 i_1867 (.ZN (n_327), .A1 (inputB[28]), .A2 (inputA[20]));
XNOR2_X1 i_1866 (.ZN (n_319), .A (n_328), .B (n_327));
AOI22_X1 i_1865 (.ZN (n_318), .A1 (n_381), .A2 (n_376), .B1 (n_375), .B2 (n_359));
AOI21_X1 i_1864 (.ZN (n_317), .A (n_333), .B1 (n_331), .B2 (n_319));
NAND2_X1 i_1863 (.ZN (n_316), .A1 (n_318), .A2 (n_317));
OAI21_X1 i_1862 (.ZN (n_315), .A (n_316), .B1 (n_318), .B2 (n_317));
INV_X1 i_1861 (.ZN (n_314), .A (inputB[19]));
NOR2_X1 i_1860 (.ZN (n_313), .A1 (n_314), .A2 (n_123));
NAND2_X1 i_1859 (.ZN (n_312), .A1 (inputB[17]), .A2 (inputA[31]));
XOR2_X1 i_1858 (.Z (n_311), .A (n_313), .B (n_312));
NAND2_X1 i_1857 (.ZN (n_310), .A1 (inputB[18]), .A2 (inputA[30]));
INV_X1 i_1856 (.ZN (n_309), .A (n_310));
AOI22_X1 i_1855 (.ZN (n_308), .A1 (n_313), .A2 (n_312), .B1 (n_311), .B2 (n_309));
NAND2_X1 i_1854 (.ZN (n_307), .A1 (inputB[18]), .A2 (inputA[31]));
XOR2_X1 i_1853 (.Z (n_305), .A (n_308), .B (n_307));
INV_X1 i_1852 (.ZN (n_304), .A (n_305));
NOR2_X1 i_1851 (.ZN (n_303), .A1 (n_314), .A2 (n_124));
XOR2_X1 i_1850 (.Z (n_302), .A (n_305), .B (n_303));
NAND2_X1 i_1849 (.ZN (n_301), .A1 (inputB[21]), .A2 (inputA[26]));
NAND2_X1 i_1848 (.ZN (n_300), .A1 (inputB[20]), .A2 (inputA[27]));
XNOR2_X1 i_1847 (.ZN (n_287), .A (n_301), .B (n_300));
NAND2_X1 i_1846 (.ZN (n_286), .A1 (inputB[22]), .A2 (inputA[25]));
NAND2_X1 i_1845 (.ZN (n_285), .A1 (inputB[17]), .A2 (inputA[29]));
NOR2_X1 i_1844 (.ZN (n_284), .A1 (n_310), .A2 (n_285));
AOI22_X1 i_1843 (.ZN (n_283), .A1 (inputB[18]), .A2 (inputA[29]), .B1 (inputB[17]), .B2 (inputA[30]));
NOR2_X1 i_1842 (.ZN (n_282), .A1 (n_284), .A2 (n_283));
NOR2_X1 i_1841 (.ZN (n_281), .A1 (n_314), .A2 (n_122));
AOI21_X1 i_1840 (.ZN (n_280), .A (n_284), .B1 (n_282), .B2 (n_281));
INV_X1 i_1839 (.ZN (n_279), .A (n_280));
OAI22_X1 i_1838 (.ZN (n_278), .A1 (n_301), .A2 (n_300), .B1 (n_287), .B2 (n_286));
XOR2_X1 i_1837 (.Z (n_277), .A (n_279), .B (n_278));
NAND2_X1 i_1836 (.ZN (n_276), .A1 (inputB[23]), .A2 (inputA[23]));
NAND2_X1 i_1835 (.ZN (n_275), .A1 (inputB[24]), .A2 (inputA[24]));
AOI22_X1 i_1834 (.ZN (n_274), .A1 (inputB[23]), .A2 (inputA[24]), .B1 (inputB[24]), .B2 (inputA[23]));
INV_X1 i_1833 (.ZN (n_273), .A (n_274));
OAI21_X1 i_1832 (.ZN (n_272), .A (n_273), .B1 (n_276), .B2 (n_275));
NAND2_X1 i_1830 (.ZN (n_271), .A1 (inputB[25]), .A2 (inputA[22]));
OAI22_X1 i_1829 (.ZN (n_270), .A1 (n_276), .A2 (n_275), .B1 (n_272), .B2 (n_271));
AOI22_X1 i_1828 (.ZN (n_269), .A1 (n_279), .A2 (n_278), .B1 (n_277), .B2 (n_270));
NAND2_X1 i_1827 (.ZN (n_268), .A1 (inputB[29]), .A2 (inputA[18]));
NAND2_X1 i_1826 (.ZN (n_267), .A1 (inputB[30]), .A2 (inputA[19]));
NOR2_X1 i_1825 (.ZN (n_266), .A1 (n_268), .A2 (n_267));
AOI22_X1 i_1824 (.ZN (n_265), .A1 (inputB[30]), .A2 (inputA[18]), .B1 (inputB[29]), .B2 (inputA[19]));
NOR2_X1 i_1823 (.ZN (n_264), .A1 (n_266), .A2 (n_265));
NAND2_X1 i_1822 (.ZN (n_263), .A1 (inputB[31]), .A2 (inputA[17]));
AOI21_X1 i_1821 (.ZN (n_262), .A (n_266), .B1 (n_264), .B2 (n_263));
XOR2_X1 i_1820 (.Z (n_261), .A (n_269), .B (n_262));
XOR2_X1 i_1819 (.Z (n_260), .A (n_302), .B (n_261));
INV_X1 i_1818 (.ZN (n_259), .A (inputA[22]));
AOI22_X1 i_1817 (.ZN (n_258), .A1 (inputB[23]), .A2 (inputA[27]), .B1 (inputB[24]), .B2 (inputA[26]));
NOR2_X1 i_1816 (.ZN (n_257), .A1 (n_218), .A2 (n_214));
NAND3_X1 i_1815 (.ZN (n_256), .A1 (inputB[24]), .A2 (n_257), .A3 (inputA[27]));
NAND2_X1 i_1814 (.ZN (n_255), .A1 (inputB[25]), .A2 (inputA[25]));
AOI22_X1 i_1813 (.ZN (n_254), .A1 (inputB[21]), .A2 (inputA[29]), .B1 (inputB[20]), .B2 (inputA[30]));
NAND3_X1 i_1812 (.ZN (n_246), .A1 (inputB[20]), .A2 (n_212), .A3 (inputA[29]));
NAND2_X1 i_1811 (.ZN (n_239), .A1 (inputB[22]), .A2 (inputA[28]));
AOI21_X1 i_1810 (.ZN (n_238), .A (n_258), .B1 (n_256), .B2 (n_255));
AOI21_X1 i_1809 (.ZN (n_237), .A (n_254), .B1 (n_246), .B2 (n_239));
NAND2_X1 i_1808 (.ZN (n_230), .A1 (n_238), .A2 (n_237));
OAI21_X1 i_1807 (.ZN (n_228), .A (n_230), .B1 (n_238), .B2 (n_237));
NAND2_X1 i_1806 (.ZN (n_227), .A1 (inputB[27]), .A2 (inputA[23]));
NOR2_X1 i_1805 (.ZN (n_226), .A1 (n_184), .A2 (n_227));
AOI21_X1 i_1804 (.ZN (n_225), .A (n_226), .B1 (n_184), .B2 (n_227));
NOR2_X1 i_1803 (.ZN (n_224), .A1 (n_259), .A2 (n_127));
AOI21_X1 i_1802 (.ZN (n_223), .A (n_226), .B1 (n_225), .B2 (n_224));
OAI21_X1 i_1801 (.ZN (n_222), .A (n_230), .B1 (n_228), .B2 (n_223));
INV_X1 i_1800 (.ZN (n_221), .A (n_222));
INV_X1 i_1799 (.ZN (n_219), .A (inputB[25]));
INV_X1 i_1798 (.ZN (n_218), .A (inputB[23]));
INV_X1 i_1797 (.ZN (n_217), .A (inputB[22]));
INV_X1 i_1796 (.ZN (n_216), .A (inputB[21]));
INV_X1 i_1795 (.ZN (n_215), .A (inputA[27]));
INV_X1 i_1794 (.ZN (n_214), .A (inputA[26]));
INV_X1 i_1793 (.ZN (n_213), .A (inputA[23]));
NOR2_X1 i_1792 (.ZN (n_212), .A1 (n_216), .A2 (n_124));
NAND2_X1 i_1791 (.ZN (n_211), .A1 (inputB[20]), .A2 (inputA[31]));
XOR2_X1 i_1790 (.Z (n_210), .A (n_212), .B (n_211));
NOR2_X1 i_1789 (.ZN (n_209), .A1 (n_217), .A2 (n_123));
NAND2_X1 i_1788 (.ZN (n_208), .A1 (inputB[21]), .A2 (inputA[31]));
AOI22_X1 i_1787 (.ZN (n_207), .A1 (n_212), .A2 (n_211), .B1 (n_210), .B2 (n_209));
INV_X1 i_1786 (.ZN (n_206), .A (n_207));
XOR2_X1 i_1785 (.Z (n_205), .A (n_208), .B (n_206));
NOR2_X1 i_1784 (.ZN (n_204), .A1 (n_217), .A2 (n_124));
NAND2_X1 i_1783 (.ZN (n_203), .A1 (inputB[29]), .A2 (inputA[23]));
INV_X1 i_1782 (.ZN (n_202), .A (n_203));
NAND2_X1 i_1781 (.ZN (n_201), .A1 (inputB[31]), .A2 (inputA[21]));
NOR2_X1 i_1780 (.ZN (n_200), .A1 (n_202), .A2 (n_201));
AOI21_X1 i_1779 (.ZN (n_196), .A (n_200), .B1 (n_202), .B2 (n_201));
NAND2_X1 i_1778 (.ZN (n_195), .A1 (inputB[30]), .A2 (inputA[22]));
INV_X1 i_1777 (.ZN (n_194), .A (n_195));
AOI22_X1 i_1776 (.ZN (n_193), .A1 (n_208), .A2 (n_206), .B1 (n_205), .B2 (n_204));
AOI22_X1 i_1775 (.ZN (n_192), .A1 (n_202), .A2 (n_201), .B1 (n_196), .B2 (n_194));
NOR2_X1 i_1774 (.ZN (n_191), .A1 (n_193), .A2 (n_192));
AOI21_X1 i_1773 (.ZN (n_190), .A (n_191), .B1 (n_193), .B2 (n_192));
NAND2_X1 i_1772 (.ZN (n_189), .A1 (inputB[24]), .A2 (inputA[28]));
AND2_X1 i_1771 (.ZN (n_188), .A1 (inputB[23]), .A2 (inputA[28]));
AND2_X1 i_1770 (.ZN (n_187), .A1 (inputB[24]), .A2 (inputA[27]));
XOR2_X1 i_1769 (.Z (n_186), .A (n_188), .B (n_187));
NOR2_X1 i_1768 (.ZN (n_185), .A1 (n_219), .A2 (n_214));
NAND2_X1 i_1767 (.ZN (n_184), .A1 (inputB[26]), .A2 (inputA[24]));
NAND2_X1 i_1766 (.ZN (n_183), .A1 (inputB[27]), .A2 (inputA[25]));
NOR2_X1 i_1765 (.ZN (n_182), .A1 (n_184), .A2 (n_183));
AOI22_X1 i_1764 (.ZN (n_181), .A1 (inputB[26]), .A2 (inputA[25]), .B1 (inputB[27]), .B2 (inputA[24]));
NOR2_X1 i_1763 (.ZN (n_180), .A1 (n_182), .A2 (n_181));
NOR2_X1 i_1762 (.ZN (n_179), .A1 (n_213), .A2 (n_127));
AOI21_X1 i_1761 (.ZN (n_178), .A (n_182), .B1 (n_180), .B2 (n_179));
AOI22_X1 i_1760 (.ZN (n_177), .A1 (n_188), .A2 (n_187), .B1 (n_186), .B2 (n_185));
XNOR2_X1 i_1759 (.ZN (n_176), .A (n_178), .B (n_177));
NAND2_X1 i_1758 (.ZN (n_175), .A1 (inputB[29]), .A2 (inputA[21]));
NOR2_X1 i_1757 (.ZN (n_174), .A1 (n_195), .A2 (n_175));
AOI22_X1 i_1756 (.ZN (n_173), .A1 (inputB[30]), .A2 (inputA[21]), .B1 (inputB[29]), .B2 (inputA[22]));
NOR2_X1 i_1755 (.ZN (n_172), .A1 (n_174), .A2 (n_173));
NAND2_X1 i_1754 (.ZN (n_171), .A1 (inputB[31]), .A2 (inputA[20]));
AOI21_X1 i_1753 (.ZN (n_170), .A (n_174), .B1 (n_172), .B2 (n_171));
OAI22_X1 i_1752 (.ZN (n_169), .A1 (n_178), .A2 (n_177), .B1 (n_176), .B2 (n_170));
AOI21_X1 i_1751 (.ZN (n_168), .A (n_191), .B1 (n_190), .B2 (n_169));
NAND2_X1 i_1750 (.ZN (n_167), .A1 (inputB[26]), .A2 (inputA[26]));
NAND2_X1 i_1749 (.ZN (n_165), .A1 (inputB[27]), .A2 (inputA[27]));
AOI22_X1 i_1748 (.ZN (n_164), .A1 (inputB[26]), .A2 (inputA[27]), .B1 (inputB[27]), .B2 (inputA[26]));
INV_X1 i_1747 (.ZN (n_158), .A (n_164));
OAI21_X1 i_1746 (.ZN (n_157), .A (n_158), .B1 (n_167), .B2 (n_165));
NAND2_X1 i_1745 (.ZN (n_156), .A1 (inputB[28]), .A2 (inputA[25]));
NAND2_X1 i_1744 (.ZN (n_155), .A1 (inputB[23]), .A2 (inputA[29]));
NAND2_X1 i_1743 (.ZN (n_154), .A1 (inputB[24]), .A2 (inputA[30]));
AOI22_X1 i_1742 (.ZN (n_153), .A1 (inputB[24]), .A2 (inputA[29]), .B1 (inputB[23]), .B2 (inputA[30]));
INV_X1 i_1741 (.ZN (n_152), .A (n_153));
OAI21_X1 i_1740 (.ZN (n_151), .A (n_152), .B1 (n_155), .B2 (n_154));
NAND2_X1 i_1739 (.ZN (n_150), .A1 (inputB[25]), .A2 (inputA[28]));
OAI22_X1 i_1738 (.ZN (n_149), .A1 (n_167), .A2 (n_165), .B1 (n_157), .B2 (n_156));
OAI22_X1 i_1737 (.ZN (n_148), .A1 (n_155), .A2 (n_154), .B1 (n_151), .B2 (n_150));
NAND2_X1 i_1736 (.ZN (n_147), .A1 (n_149), .A2 (n_148));
OAI21_X1 i_1735 (.ZN (n_146), .A (n_147), .B1 (n_149), .B2 (n_148));
NAND2_X1 i_1734 (.ZN (n_145), .A1 (inputB[30]), .A2 (inputA[24]));
NOR2_X1 i_1733 (.ZN (n_144), .A1 (n_203), .A2 (n_145));
AOI22_X1 i_1732 (.ZN (n_143), .A1 (inputB[29]), .A2 (inputA[24]), .B1 (inputB[30]), .B2 (inputA[23]));
NOR2_X1 i_1731 (.ZN (n_142), .A1 (n_144), .A2 (n_143));
NAND2_X1 i_1730 (.ZN (n_141), .A1 (inputB[31]), .A2 (inputA[22]));
AOI21_X1 i_1729 (.ZN (n_140), .A (n_144), .B1 (n_142), .B2 (n_141));
NAND2_X1 i_1728 (.ZN (n_139), .A1 (inputB[29]), .A2 (inputA[25]));
XNOR2_X1 i_1727 (.ZN (n_138), .A (n_145), .B (n_139));
NOR2_X1 i_1726 (.ZN (n_137), .A1 (n_213), .A2 (n_129));
XNOR2_X1 i_1725 (.ZN (n_136), .A (n_146), .B (n_140));
XNOR2_X1 i_1724 (.ZN (n_135), .A (n_138), .B (n_137));
NAND2_X1 i_1723 (.ZN (n_133), .A1 (n_136), .A2 (n_135));
NOR2_X1 i_1722 (.ZN (n_132), .A1 (n_136), .A2 (n_135));
AOI21_X1 i_1721 (.ZN (n_131), .A (n_132), .B1 (n_136), .B2 (n_135));
XNOR2_X1 i_1720 (.ZN (n_130), .A (n_168), .B (n_131));
INV_X1 i_1719 (.ZN (n_129), .A (inputB[31]));
INV_X1 i_1718 (.ZN (n_128), .A (inputB[29]));
INV_X1 i_1717 (.ZN (n_127), .A (inputB[28]));
INV_X1 i_1716 (.ZN (n_126), .A (inputB[27]));
INV_X1 i_1715 (.ZN (n_125), .A (inputA[31]));
INV_X1 i_1714 (.ZN (n_124), .A (inputA[30]));
INV_X1 i_1713 (.ZN (n_123), .A (inputA[29]));
INV_X1 i_1712 (.ZN (n_122), .A (inputA[28]));
NOR2_X1 i_1711 (.ZN (n_118), .A1 (n_127), .A2 (n_123));
NAND2_X1 i_1710 (.ZN (n_117), .A1 (inputB[26]), .A2 (inputA[31]));
XOR2_X1 i_1709 (.Z (n_116), .A (n_118), .B (n_117));
NOR2_X1 i_1708 (.ZN (n_115), .A1 (n_126), .A2 (n_124));
INV_X1 i_1707 (.ZN (n_114), .A (n_115));
NOR2_X1 i_1706 (.ZN (n_113), .A1 (n_126), .A2 (n_125));
AOI22_X1 i_1705 (.ZN (n_112), .A1 (n_118), .A2 (n_117), .B1 (n_116), .B2 (n_115));
NOR2_X1 i_1704 (.ZN (n_111), .A1 (n_113), .A2 (n_112));
AOI21_X1 i_1703 (.ZN (n_110), .A (n_111), .B1 (n_113), .B2 (n_112));
NOR2_X1 i_1702 (.ZN (n_109), .A1 (n_127), .A2 (n_124));
AOI21_X1 i_1701 (.ZN (n_107), .A (n_111), .B1 (n_110), .B2 (n_109));
NAND2_X1 i_1700 (.ZN (n_106), .A1 (inputB[29]), .A2 (inputA[28]));
NAND2_X1 i_1699 (.ZN (n_105), .A1 (inputB[30]), .A2 (inputA[29]));
NOR2_X1 i_1698 (.ZN (n_104), .A1 (n_106), .A2 (n_105));
AOI22_X1 i_1697 (.ZN (n_103), .A1 (inputB[29]), .A2 (inputA[29]), .B1 (inputB[30]), .B2 (inputA[28]));
NOR2_X1 i_1696 (.ZN (n_102), .A1 (n_104), .A2 (n_103));
NAND2_X1 i_1695 (.ZN (n_101), .A1 (inputB[31]), .A2 (inputA[27]));
AOI21_X1 i_1694 (.ZN (n_100), .A (n_104), .B1 (n_102), .B2 (n_101));
NOR2_X1 i_1693 (.ZN (n_99), .A1 (n_127), .A2 (n_125));
NOR2_X1 i_1692 (.ZN (n_98), .A1 (n_100), .A2 (n_99));
INV_X1 i_1691 (.ZN (n_97), .A (n_98));
AOI21_X1 i_1690 (.ZN (n_96), .A (n_98), .B1 (n_100), .B2 (n_99));
AOI22_X1 i_1689 (.ZN (n_92), .A1 (n_100), .A2 (n_99), .B1 (n_107), .B2 (n_97));
NAND2_X1 i_1688 (.ZN (n_91), .A1 (inputB[30]), .A2 (inputA[30]));
NAND4_X1 i_1687 (.ZN (n_89), .A1 (inputB[29]), .A2 (inputA[29]), .A3 (inputB[30]), .A4 (inputA[30]));
OAI21_X1 i_1686 (.ZN (n_88), .A (n_105), .B1 (n_128), .B2 (n_124));
NAND2_X1 i_1685 (.ZN (n_87), .A1 (n_89), .A2 (n_88));
NOR2_X1 i_1684 (.ZN (n_86), .A1 (n_129), .A2 (n_122));
OAI21_X1 i_1683 (.ZN (n_85), .A (n_89), .B1 (n_87), .B2 (n_86));
NOR2_X1 i_1682 (.ZN (n_84), .A1 (n_128), .A2 (n_125));
XOR2_X1 i_1681 (.Z (n_83), .A (n_91), .B (n_84));
NOR2_X1 i_1680 (.ZN (n_82), .A1 (n_129), .A2 (n_123));
XNOR2_X1 i_1679 (.ZN (n_81), .A (n_83), .B (n_82));
NAND3_X1 i_1678 (.ZN (n_80), .A1 (n_92), .A2 (n_85), .A3 (n_81));
INV_X1 i_1677 (.ZN (n_79), .A (n_80));
XNOR2_X1 i_1676 (.ZN (result[3]), .A (n_74), .B (n_78));
XOR2_X1 i_1675 (.Z (n_78), .A (n_76), .B (n_77));
NAND2_X1 i_1674 (.ZN (n_77), .A1 (inputB[3]), .A2 (inputA[0]));
XNOR2_X1 i_1673 (.ZN (n_76), .A (n_75), .B (n_61));
NAND2_X1 i_1672 (.ZN (n_75), .A1 (inputB[1]), .A2 (inputA[2]));
NAND2_X1 i_1671 (.ZN (n_74), .A1 (n_72), .A2 (n_73));
NAND2_X1 i_1670 (.ZN (n_73), .A1 (n_69), .A2 (n_71));
OR2_X1 i_1669 (.ZN (n_72), .A1 (n_69), .A2 (n_71));
OAI21_X1 i_1668 (.ZN (n_71), .A (n_54), .B1 (n_70), .B2 (n_51));
INV_X1 i_1667 (.ZN (n_70), .A (n_53));
XNOR2_X1 i_1666 (.ZN (n_69), .A (n_68), .B (n_58));
NAND2_X1 i_1665 (.ZN (n_68), .A1 (inputB[0]), .A2 (inputA[3]));
INV_X1 i_1664 (.ZN (n_67), .A (inputA[2]));
INV_X1 i_1663 (.ZN (n_66), .A (inputA[0]));
INV_X1 i_1662 (.ZN (n_63), .A (inputB[1]));
INV_X1 i_1661 (.ZN (n_62), .A (inputB[0]));
NAND2_X1 i_1660 (.ZN (n_61), .A1 (inputA[1]), .A2 (inputB[2]));
AND2_X1 i_1659 (.ZN (n_60), .A1 (inputA[0]), .A2 (inputB[2]));
AND2_X1 i_1658 (.ZN (n_59), .A1 (inputA[1]), .A2 (inputB[1]));
NAND2_X1 i_1657 (.ZN (n_58), .A1 (n_60), .A2 (n_59));
OAI21_X1 i_1656 (.ZN (n_57), .A (n_58), .B1 (n_60), .B2 (n_59));
NAND2_X1 i_1655 (.ZN (n_56), .A1 (inputA[2]), .A2 (inputB[0]));
NAND2_X1 i_1654 (.ZN (n_54), .A1 (n_57), .A2 (n_56));
OR2_X1 i_1653 (.ZN (n_53), .A1 (n_57), .A2 (n_56));
NAND2_X1 i_1652 (.ZN (n_52), .A1 (n_54), .A2 (n_53));
NOR2_X1 i_1651 (.ZN (result[0]), .A1 (n_66), .A2 (n_62));
AND2_X1 i_1650 (.ZN (n_51), .A1 (n_59), .A2 (result[0]));
XNOR2_X1 i_1649 (.ZN (result[2]), .A (n_52), .B (n_51));
OAI21_X1 i_4711 (.ZN (result[63]), .A (n_6), .B1 (n_5), .B2 (n_8));
XNOR2_X1 i_4710 (.ZN (result[62]), .A (n_5), .B (n_8));
OAI21_X1 i_1648 (.ZN (n_8), .A (n_6), .B1 (n_4620), .B2 (n_7));
NAND3_X1 i_1647 (.ZN (n_7), .A1 (n_91), .A2 (inputB[31]), .A3 (inputA[31]));
OAI21_X1 i_1646 (.ZN (n_6), .A (n_4620), .B1 (n_129), .B2 (n_125));
NAND3_X1 i_1645 (.ZN (n_5), .A1 (n_2), .A2 (n_4), .A3 (n_0));
OAI211_X1 i_1644 (.ZN (n_4), .A (n_4610), .B (n_4627), .C1 (n_79), .C2 (n_4618));
OAI21_X1 i_1643 (.ZN (n_2), .A (n_4618), .B1 (n_4609), .B2 (n_4626));
XNOR2_X1 i_4703 (.ZN (result[61]), .A (n_1), .B (n_4618));
OAI211_X1 i_4694 (.ZN (n_1), .A (n_4631), .B (n_0), .C1 (n_4609), .C2 (n_4627));
NAND2_X1 i_1642 (.ZN (n_0), .A1 (n_4609), .A2 (n_4626));
AOI22_X1 i_4692 (.ZN (n_4631), .A1 (n_4611), .A2 (n_4625), .B1 (n_4610), .B2 (n_79));
XOR2_X1 i_4690 (.Z (result[60]), .A (n_4612), .B (n_4629));
OAI21_X1 i_4689 (.ZN (n_4629), .A (n_80), .B1 (n_4626), .B2 (n_4628));
INV_X1 i_4688 (.ZN (n_4628), .A (n_4627));
OR2_X1 i_1641 (.ZN (n_4627), .A1 (n_92), .A2 (n_4624));
INV_X1 i_1640 (.ZN (n_4626), .A (n_4625));
AOI22_X1 i_1639 (.ZN (n_4625), .A1 (n_92), .A2 (n_4624), .B1 (n_81), .B2 (n_85));
OR2_X1 i_1638 (.ZN (n_4624), .A1 (n_81), .A2 (n_85));
NOR2_X1 i_4672 (.ZN (n_4612), .A1 (n_4609), .A2 (n_4611));
INV_X1 i_4671 (.ZN (n_4611), .A (n_4610));
NAND2_X1 i_1637 (.ZN (n_4610), .A1 (n_4607), .A2 (n_4608));
NOR2_X1 i_1636 (.ZN (n_4609), .A1 (n_4607), .A2 (n_4608));
OAI22_X1 i_1635 (.ZN (n_4608), .A1 (n_4603), .A2 (n_4604), .B1 (n_4598), .B2 (n_4602));
OAI22_X1 i_1634 (.ZN (n_4607), .A1 (n_4591), .A2 (n_4606), .B1 (n_4592), .B2 (n_4605));
XNOR2_X1 i_4666 (.ZN (result[59]), .A (n_4591), .B (n_4606));
XNOR2_X1 i_1633 (.ZN (n_4606), .A (n_4592), .B (n_4605));
XNOR2_X1 i_1632 (.ZN (n_4605), .A (n_4603), .B (n_4604));
AOI22_X1 i_1631 (.ZN (n_4604), .A1 (n_4570), .A2 (n_4579), .B1 (n_4576), .B2 (n_4578));
XNOR2_X1 i_1630 (.ZN (n_4603), .A (n_4598), .B (n_4602));
XOR2_X1 i_1629 (.Z (n_4602), .A (n_87), .B (n_86));
XNOR2_X1 i_1628 (.ZN (n_4598), .A (n_107), .B (n_96));
AOI22_X1 i_1627 (.ZN (n_4592), .A1 (n_4585), .A2 (n_4584), .B1 (n_4583), .B2 (n_4580));
AOI21_X1 i_1626 (.ZN (n_4591), .A (n_4589), .B1 (n_4561), .B2 (n_4587));
XNOR2_X1 i_4649 (.ZN (result[58]), .A (n_4561), .B (n_4590));
NOR2_X1 i_4648 (.ZN (n_4590), .A1 (n_4588), .A2 (n_4589));
NOR2_X1 i_1625 (.ZN (n_4589), .A1 (n_4617), .A2 (n_4586));
INV_X1 i_4646 (.ZN (n_4588), .A (n_4587));
NAND2_X1 i_1624 (.ZN (n_4587), .A1 (n_4617), .A2 (n_4586));
XNOR2_X1 i_1623 (.ZN (n_4586), .A (n_4584), .B (n_4585));
AOI22_X1 i_1622 (.ZN (n_4585), .A1 (n_4597), .A2 (n_4615), .B1 (n_4599), .B2 (n_4614));
XOR2_X1 i_1621 (.Z (n_4584), .A (n_4580), .B (n_4583));
AOI22_X1 i_1620 (.ZN (n_4583), .A1 (n_4581), .A2 (n_4596), .B1 (n_4594), .B2 (n_4582));
INV_X1 i_1619 (.ZN (n_4582), .A (n_4595));
INV_X1 i_1618 (.ZN (n_4581), .A (n_4593));
XOR2_X1 i_1617 (.Z (n_4580), .A (n_4570), .B (n_4579));
XOR2_X1 i_1616 (.Z (n_4579), .A (n_4576), .B (n_4578));
AOI22_X1 i_1615 (.ZN (n_4578), .A1 (n_4601), .A2 (n_4613), .B1 (n_4577), .B2 (n_4600));
INV_X1 i_1614 (.ZN (n_4577), .A (n_106));
XNOR2_X1 i_1613 (.ZN (n_4576), .A (n_102), .B (n_101));
XNOR2_X1 i_1612 (.ZN (n_4570), .A (n_110), .B (n_109));
OAI21_X1 i_1611 (.ZN (n_4561), .A (n_4559), .B1 (n_4537), .B2 (n_4560));
XNOR2_X1 i_4618 (.ZN (result[57]), .A (n_4537), .B (n_4560));
OAI21_X1 i_1610 (.ZN (n_4560), .A (n_4559), .B1 (n_4538), .B2 (n_4558));
NAND2_X1 i_1609 (.ZN (n_4559), .A1 (n_4538), .A2 (n_4558));
XNOR2_X1 i_1608 (.ZN (n_4558), .A (n_4575), .B (n_4616));
AOI22_X1 i_1607 (.ZN (n_4538), .A1 (n_4524), .A2 (n_4533), .B1 (n_4481), .B2 (n_4521));
AOI22_X1 i_1606 (.ZN (n_4537), .A1 (n_4505), .A2 (n_4535), .B1 (n_4536), .B2 (n_4534));
INV_X1 i_1605 (.ZN (n_4536), .A (n_4506));
XNOR2_X1 i_4592 (.ZN (result[56]), .A (n_4505), .B (n_4535));
XNOR2_X1 i_1604 (.ZN (n_4535), .A (n_4506), .B (n_4534));
XNOR2_X1 i_1603 (.ZN (n_4534), .A (n_4524), .B (n_4533));
XNOR2_X1 i_1602 (.ZN (n_4533), .A (n_4532), .B (n_4552));
XOR2_X1 i_1601 (.Z (n_4524), .A (n_4521), .B (n_4481));
XOR2_X1 i_1600 (.Z (n_4521), .A (n_4565), .B (n_4571));
AOI22_X1 i_1599 (.ZN (n_4506), .A1 (n_4499), .A2 (n_4500), .B1 (n_4479), .B2 (n_4498));
AOI22_X1 i_1598 (.ZN (n_4505), .A1 (n_4469), .A2 (n_4504), .B1 (n_4503), .B2 (n_4501));
XOR2_X1 i_4560 (.Z (result[55]), .A (n_4469), .B (n_4504));
XOR2_X1 i_1597 (.Z (n_4504), .A (n_4501), .B (n_4503));
AOI22_X1 i_1596 (.ZN (n_4503), .A1 (n_4463), .A2 (n_4502), .B1 (n_4461), .B2 (n_4462));
INV_X1 i_1595 (.ZN (n_4502), .A (n_4465));
XNOR2_X1 i_1594 (.ZN (n_4501), .A (n_4499), .B (n_4500));
AOI22_X1 i_1593 (.ZN (n_4500), .A1 (n_4442), .A2 (n_130), .B1 (n_4440), .B2 (n_4441));
XOR2_X1 i_1592 (.Z (n_4499), .A (n_4479), .B (n_4498));
XNOR2_X1 i_1591 (.ZN (n_4498), .A (n_4549), .B (n_4551));
XOR2_X1 i_1590 (.Z (n_4479), .A (n_4483), .B (n_4482));
AOI22_X1 i_1589 (.ZN (n_4469), .A1 (n_4429), .A2 (n_4468), .B1 (n_4466), .B2 (n_4467));
XNOR2_X1 i_4523 (.ZN (result[54]), .A (n_4429), .B (n_4468));
XOR2_X1 i_1588 (.Z (n_4468), .A (n_4466), .B (n_4467));
AOI22_X1 i_1587 (.ZN (n_4467), .A1 (n_4425), .A2 (n_4426), .B1 (n_4424), .B2 (n_4398));
XNOR2_X1 i_1586 (.ZN (n_4466), .A (n_4463), .B (n_4465));
AOI22_X1 i_1585 (.ZN (n_4465), .A1 (n_4400), .A2 (n_4423), .B1 (n_4464), .B2 (n_4422));
INV_X1 i_1584 (.ZN (n_4464), .A (n_4401));
XOR2_X1 i_1583 (.Z (n_4463), .A (n_4461), .B (n_4462));
OAI21_X1 i_1582 (.ZN (n_4462), .A (n_4394), .B1 (n_4395), .B2 (n_4397));
XNOR2_X1 i_1581 (.ZN (n_4461), .A (n_4442), .B (n_130));
XOR2_X1 i_1580 (.Z (n_4442), .A (n_4440), .B (n_4441));
OAI21_X1 i_1579 (.ZN (n_4441), .A (n_4414), .B1 (n_4415), .B2 (n_4421));
XNOR2_X1 i_1578 (.ZN (n_4440), .A (n_4496), .B (n_4491));
OAI22_X1 i_1577 (.ZN (n_4429), .A1 (n_4378), .A2 (n_4427), .B1 (n_4377), .B2 (n_4428));
INV_X1 i_1576 (.ZN (n_4428), .A (n_4375));
XNOR2_X1 i_4481 (.ZN (result[53]), .A (n_4378), .B (n_4427));
XOR2_X1 i_1575 (.Z (n_4427), .A (n_4425), .B (n_4426));
AOI22_X1 i_1574 (.ZN (n_4426), .A1 (n_4360), .A2 (n_4359), .B1 (n_4343), .B2 (n_4358));
XOR2_X1 i_1573 (.Z (n_4425), .A (n_4398), .B (n_4424));
XNOR2_X1 i_1572 (.ZN (n_4424), .A (n_4400), .B (n_4423));
XNOR2_X1 i_1571 (.ZN (n_4423), .A (n_4401), .B (n_4422));
XNOR2_X1 i_1570 (.ZN (n_4422), .A (n_4415), .B (n_4421));
XNOR2_X1 i_1569 (.ZN (n_4421), .A (n_157), .B (n_156));
OAI21_X1 i_1568 (.ZN (n_4415), .A (n_4414), .B1 (n_4407), .B2 (n_4413));
NAND2_X1 i_1567 (.ZN (n_4414), .A1 (n_4407), .A2 (n_4413));
XOR2_X1 i_1566 (.Z (n_4413), .A (n_142), .B (n_141));
XOR2_X1 i_1565 (.Z (n_4407), .A (n_151), .B (n_150));
AOI22_X1 i_1564 (.ZN (n_4401), .A1 (n_4348), .A2 (n_4357), .B1 (n_4352), .B2 (n_4356));
OAI22_X1 i_1563 (.ZN (n_4400), .A1 (n_4447), .A2 (n_4420), .B1 (n_4399), .B2 (n_4430));
INV_X1 i_1562 (.ZN (n_4399), .A (n_4438));
XNOR2_X1 i_1561 (.ZN (n_4398), .A (n_4395), .B (n_4397));
OAI22_X1 i_1560 (.ZN (n_4397), .A1 (n_4341), .A2 (n_221), .B1 (n_4336), .B2 (n_4340));
OAI21_X1 i_1559 (.ZN (n_4395), .A (n_4394), .B1 (n_4383), .B2 (n_4393));
NAND2_X1 i_1558 (.ZN (n_4394), .A1 (n_4383), .A2 (n_4393));
XNOR2_X1 i_1557 (.ZN (n_4393), .A (n_190), .B (n_169));
XNOR2_X1 i_1556 (.ZN (n_4383), .A (n_4513), .B (n_4511));
XOR2_X1 i_1555 (.Z (n_4378), .A (n_4375), .B (n_4377));
OAI22_X1 i_1554 (.ZN (n_4377), .A1 (n_4331), .A2 (n_4374), .B1 (n_4376), .B2 (n_4372));
INV_X1 i_1553 (.ZN (n_4376), .A (n_4373));
OAI21_X1 i_1552 (.ZN (n_4375), .A (n_4370), .B1 (n_4371), .B2 (n_4361));
XOR2_X1 i_4427 (.Z (result[52]), .A (n_4331), .B (n_4374));
XOR2_X1 i_1551 (.Z (n_4374), .A (n_4372), .B (n_4373));
OAI21_X1 i_1550 (.ZN (n_4373), .A (n_4323), .B1 (n_4326), .B2 (n_4324));
XOR2_X1 i_1549 (.Z (n_4372), .A (n_4361), .B (n_4371));
OAI21_X1 i_1548 (.ZN (n_4371), .A (n_4370), .B1 (n_4363), .B2 (n_4419));
NAND2_X1 i_1547 (.ZN (n_4370), .A1 (n_4363), .A2 (n_4419));
AOI22_X1 i_1546 (.ZN (n_4363), .A1 (n_4362), .A2 (n_4305), .B1 (n_4283), .B2 (n_4304));
INV_X1 i_1545 (.ZN (n_4362), .A (n_4270));
XNOR2_X1 i_1544 (.ZN (n_4361), .A (n_4359), .B (n_4360));
AOI22_X1 i_1543 (.ZN (n_4360), .A1 (n_4318), .A2 (n_4380), .B1 (n_4307), .B2 (n_4317));
XOR2_X1 i_1542 (.Z (n_4359), .A (n_4343), .B (n_4358));
XOR2_X1 i_1541 (.Z (n_4358), .A (n_4348), .B (n_4357));
XOR2_X1 i_1540 (.Z (n_4357), .A (n_4352), .B (n_4356));
XNOR2_X1 i_1539 (.ZN (n_4356), .A (n_4512), .B (n_4355));
NAND2_X1 i_1538 (.ZN (n_4355), .A1 (inputA[24]), .A2 (inputB[28]));
XOR2_X1 i_1537 (.Z (n_4352), .A (n_196), .B (n_195));
XNOR2_X1 i_1536 (.ZN (n_4348), .A (n_176), .B (n_170));
XOR2_X1 i_1535 (.Z (n_4343), .A (n_4341), .B (n_222));
XNOR2_X1 i_1534 (.ZN (n_4341), .A (n_4336), .B (n_4340));
XNOR2_X1 i_1533 (.ZN (n_4340), .A (n_4516), .B (n_4339));
NAND2_X1 i_1532 (.ZN (n_4339), .A1 (inputB[25]), .A2 (inputA[27]));
XNOR2_X1 i_1531 (.ZN (n_4336), .A (n_205), .B (n_204));
OAI22_X1 i_1530 (.ZN (n_4331), .A1 (n_4268), .A2 (n_4329), .B1 (n_4330), .B2 (n_4327));
INV_X1 i_1529 (.ZN (n_4330), .A (n_4328));
XNOR2_X1 i_4381 (.ZN (result[51]), .A (n_4268), .B (n_4329));
XOR2_X1 i_1528 (.Z (n_4329), .A (n_4327), .B (n_4328));
AOI22_X1 i_1527 (.ZN (n_4328), .A1 (n_4252), .A2 (n_4265), .B1 (n_4212), .B2 (n_4251));
XOR2_X1 i_1526 (.Z (n_4327), .A (n_4324), .B (n_4326));
AOI22_X1 i_1525 (.ZN (n_4326), .A1 (n_4325), .A2 (n_4264), .B1 (n_4263), .B2 (n_4262));
INV_X1 i_1524 (.ZN (n_4325), .A (n_4253));
OAI21_X1 i_1523 (.ZN (n_4324), .A (n_4323), .B1 (n_4306), .B2 (n_4322));
NAND2_X1 i_1522 (.ZN (n_4323), .A1 (n_4306), .A2 (n_4322));
XOR2_X1 i_1521 (.Z (n_4322), .A (n_4318), .B (n_4380));
XOR2_X1 i_1520 (.Z (n_4318), .A (n_4307), .B (n_4317));
XNOR2_X1 i_1519 (.ZN (n_4317), .A (n_4431), .B (n_4437));
AOI22_X1 i_1518 (.ZN (n_4307), .A1 (n_4219), .A2 (n_4229), .B1 (n_4228), .B2 (n_4223));
XNOR2_X1 i_1517 (.ZN (n_4306), .A (n_4270), .B (n_4305));
XOR2_X1 i_1516 (.Z (n_4305), .A (n_4283), .B (n_4304));
OAI21_X1 i_1515 (.ZN (n_4304), .A (n_4439), .B1 (n_4444), .B2 (n_4443));
XNOR2_X1 i_1514 (.ZN (n_4283), .A (n_4457), .B (n_4448));
AOI22_X1 i_1513 (.ZN (n_4270), .A1 (n_4231), .A2 (n_4250), .B1 (n_4269), .B2 (n_4230));
INV_X1 i_1512 (.ZN (n_4269), .A (n_4213));
AOI22_X1 i_1511 (.ZN (n_4268), .A1 (n_4209), .A2 (n_4267), .B1 (n_4266), .B2 (n_4210));
XNOR2_X1 i_4318 (.ZN (result[50]), .A (n_4209), .B (n_4267));
XOR2_X1 i_1510 (.Z (n_4267), .A (n_4210), .B (n_4266));
XNOR2_X1 i_1509 (.ZN (n_4266), .A (n_4252), .B (n_4265));
XNOR2_X1 i_1508 (.ZN (n_4265), .A (n_4253), .B (n_4264));
XOR2_X1 i_1507 (.Z (n_4264), .A (n_4262), .B (n_4263));
OAI21_X1 i_1506 (.ZN (n_4263), .A (n_316), .B1 (n_315), .B2 (n_260));
XOR2_X1 i_1505 (.Z (n_4262), .A (n_4384), .B (n_4382));
AOI22_X1 i_1504 (.ZN (n_4253), .A1 (n_4183), .A2 (n_4166), .B1 (n_4182), .B2 (n_415));
XOR2_X1 i_1503 (.Z (n_4252), .A (n_4212), .B (n_4251));
XOR2_X1 i_1502 (.Z (n_4251), .A (n_4231), .B (n_4250));
XNOR2_X1 i_1501 (.ZN (n_4250), .A (n_4451), .B (n_4249));
NOR2_X1 i_1500 (.ZN (n_4249), .A1 (n_4247), .A2 (n_4449));
INV_X1 i_1499 (.ZN (n_4247), .A (n_4452));
XNOR2_X1 i_1498 (.ZN (n_4231), .A (n_4213), .B (n_4230));
XNOR2_X1 i_1497 (.ZN (n_4230), .A (n_4219), .B (n_4229));
XOR2_X1 i_1496 (.Z (n_4229), .A (n_4223), .B (n_4228));
XNOR2_X1 i_1495 (.ZN (n_4228), .A (n_4435), .B (n_4434));
XNOR2_X1 i_1494 (.ZN (n_4223), .A (n_225), .B (n_224));
XNOR2_X1 i_1493 (.ZN (n_4219), .A (n_4473), .B (n_4470));
AOI22_X1 i_1492 (.ZN (n_4213), .A1 (n_426), .A2 (n_416), .B1 (n_421), .B2 (n_417));
OAI22_X1 i_1491 (.ZN (n_4212), .A1 (n_4204), .A2 (n_4202), .B1 (n_4211), .B2 (n_4201));
INV_X1 i_1490 (.ZN (n_4211), .A (n_4186));
AOI22_X1 i_1489 (.ZN (n_4210), .A1 (n_4185), .A2 (n_4205), .B1 (n_4148), .B2 (n_4184));
OAI22_X1 i_1488 (.ZN (n_4209), .A1 (n_4145), .A2 (n_4207), .B1 (n_4208), .B2 (n_4206));
INV_X1 i_1487 (.ZN (n_4208), .A (n_4146));
XNOR2_X1 i_4257 (.ZN (result[49]), .A (n_4145), .B (n_4207));
XOR2_X1 i_1486 (.Z (n_4207), .A (n_4146), .B (n_4206));
XOR2_X1 i_1485 (.Z (n_4206), .A (n_4185), .B (n_4205));
XOR2_X1 i_1484 (.Z (n_4205), .A (n_4202), .B (n_4204));
AOI22_X1 i_1483 (.ZN (n_4204), .A1 (n_4203), .A2 (n_4138), .B1 (n_4137), .B2 (n_4122));
INV_X1 i_1482 (.ZN (n_4203), .A (n_4106));
XOR2_X1 i_1481 (.Z (n_4202), .A (n_4186), .B (n_4201));
XNOR2_X1 i_1480 (.ZN (n_4201), .A (n_315), .B (n_260));
OAI21_X1 i_1479 (.ZN (n_4186), .A (n_4084), .B1 (n_4085), .B2 (n_484));
XOR2_X1 i_1478 (.Z (n_4185), .A (n_4148), .B (n_4184));
XOR2_X1 i_1477 (.Z (n_4184), .A (n_4166), .B (n_4183));
XOR2_X1 i_1476 (.Z (n_4183), .A (n_415), .B (n_4182));
AOI22_X1 i_1475 (.ZN (n_4182), .A1 (n_4101), .A2 (n_4181), .B1 (n_4092), .B2 (n_4100));
INV_X1 i_1474 (.ZN (n_4181), .A (n_4102));
XNOR2_X1 i_1473 (.ZN (n_4166), .A (n_4405), .B (n_4392));
AOI22_X1 i_1472 (.ZN (n_4148), .A1 (n_4147), .A2 (n_4104), .B1 (n_4087), .B2 (n_4103));
INV_X1 i_1471 (.ZN (n_4147), .A (n_4080));
AOI22_X1 i_1470 (.ZN (n_4146), .A1 (n_4140), .A2 (n_4141), .B1 (n_4105), .B2 (n_4139));
AOI22_X1 i_1469 (.ZN (n_4145), .A1 (n_4077), .A2 (n_4143), .B1 (n_4144), .B2 (n_4142));
INV_X1 i_1468 (.ZN (n_4144), .A (n_4079));
XNOR2_X1 i_4192 (.ZN (result[48]), .A (n_4077), .B (n_4143));
XNOR2_X1 i_1467 (.ZN (n_4143), .A (n_4079), .B (n_4142));
XNOR2_X1 i_1466 (.ZN (n_4142), .A (n_4140), .B (n_4141));
AOI22_X1 i_1465 (.ZN (n_4141), .A1 (n_4021), .A2 (n_4022), .B1 (n_4019), .B2 (n_4020));
XOR2_X1 i_1464 (.Z (n_4140), .A (n_4105), .B (n_4139));
XNOR2_X1 i_1463 (.ZN (n_4139), .A (n_4106), .B (n_4138));
XOR2_X1 i_1462 (.Z (n_4138), .A (n_4122), .B (n_4137));
XNOR2_X1 i_1461 (.ZN (n_4137), .A (n_375), .B (n_359));
XNOR2_X1 i_1460 (.ZN (n_4122), .A (n_331), .B (n_319));
AOI22_X1 i_1459 (.ZN (n_4106), .A1 (n_4017), .A2 (n_4018), .B1 (n_4016), .B2 (n_4015));
XOR2_X1 i_1458 (.Z (n_4105), .A (n_4080), .B (n_4104));
XOR2_X1 i_1457 (.Z (n_4104), .A (n_4087), .B (n_4103));
XNOR2_X1 i_1456 (.ZN (n_4103), .A (n_4101), .B (n_4102));
AOI22_X1 i_1455 (.ZN (n_4102), .A1 (n_4048), .A2 (n_4054), .B1 (n_4043), .B2 (n_4047));
XOR2_X1 i_1454 (.Z (n_4101), .A (n_4092), .B (n_4100));
XNOR2_X1 i_1453 (.ZN (n_4100), .A (n_277), .B (n_270));
XNOR2_X1 i_1452 (.ZN (n_4092), .A (n_440), .B (n_427));
XNOR2_X1 i_1451 (.ZN (n_4087), .A (n_4085), .B (n_484));
OAI21_X1 i_1450 (.ZN (n_4085), .A (n_4084), .B1 (n_531), .B2 (n_4081));
NAND2_X1 i_1449 (.ZN (n_4084), .A1 (n_4081), .A2 (n_531));
OAI22_X1 i_1448 (.ZN (n_4081), .A1 (n_4012), .A2 (n_4014), .B1 (n_4005), .B2 (n_4011));
AOI22_X1 i_1447 (.ZN (n_4080), .A1 (n_4056), .A2 (n_4068), .B1 (n_4038), .B2 (n_4055));
AOI22_X1 i_1446 (.ZN (n_4079), .A1 (n_4070), .A2 (n_4078), .B1 (n_4023), .B2 (n_4069));
INV_X1 i_1445 (.ZN (n_4078), .A (n_4072));
OAI22_X1 i_1444 (.ZN (n_4077), .A1 (n_4004), .A2 (n_4075), .B1 (n_4073), .B2 (n_4076));
INV_X1 i_1443 (.ZN (n_4076), .A (n_4074));
XNOR2_X1 i_4123 (.ZN (result[47]), .A (n_4004), .B (n_4075));
XOR2_X1 i_1442 (.Z (n_4075), .A (n_4073), .B (n_4074));
AOI22_X1 i_1441 (.ZN (n_4074), .A1 (n_4000), .A2 (n_3957), .B1 (n_3956), .B2 (n_3954));
XOR2_X1 i_1440 (.Z (n_4073), .A (n_4070), .B (n_4072));
AOI22_X1 i_1439 (.ZN (n_4072), .A1 (n_3997), .A2 (n_4071), .B1 (n_3995), .B2 (n_3996));
INV_X1 i_1438 (.ZN (n_4071), .A (n_3999));
XOR2_X1 i_1437 (.Z (n_4070), .A (n_4023), .B (n_4069));
XOR2_X1 i_1436 (.Z (n_4069), .A (n_4056), .B (n_4068));
XOR2_X1 i_1435 (.Z (n_4068), .A (n_550), .B (n_532));
XOR2_X1 i_1434 (.Z (n_4056), .A (n_4038), .B (n_4055));
XOR2_X1 i_1433 (.Z (n_4055), .A (n_4048), .B (n_4054));
XNOR2_X1 i_1432 (.ZN (n_4054), .A (n_432), .B (n_431));
XOR2_X1 i_1431 (.Z (n_4048), .A (n_4043), .B (n_4047));
XNOR2_X1 i_1430 (.ZN (n_4047), .A (n_287), .B (n_286));
XNOR2_X1 i_1429 (.ZN (n_4043), .A (n_272), .B (n_271));
XNOR2_X1 i_1428 (.ZN (n_4038), .A (n_526), .B (n_485));
XOR2_X1 i_1427 (.Z (n_4023), .A (n_4021), .B (n_4022));
AOI22_X1 i_1426 (.ZN (n_4022), .A1 (n_3931), .A2 (n_3953), .B1 (n_3925), .B2 (n_3930));
XOR2_X1 i_1425 (.Z (n_4021), .A (n_4019), .B (n_4020));
OAI21_X1 i_1424 (.ZN (n_4020), .A (n_3975), .B1 (n_3976), .B2 (n_3994));
XNOR2_X1 i_1423 (.ZN (n_4019), .A (n_4017), .B (n_4018));
OAI22_X1 i_1422 (.ZN (n_4018), .A1 (n_3929), .A2 (n_3928), .B1 (n_3926), .B2 (n_3927));
XOR2_X1 i_1421 (.Z (n_4017), .A (n_4015), .B (n_4016));
AOI22_X1 i_1420 (.ZN (n_4016), .A1 (n_3943), .A2 (n_3952), .B1 (n_3936), .B2 (n_3942));
XOR2_X1 i_1419 (.Z (n_4015), .A (n_4012), .B (n_4014));
AOI22_X1 i_1418 (.ZN (n_4014), .A1 (n_553), .A2 (n_552), .B1 (n_4013), .B2 (n_554));
INV_X1 i_1417 (.ZN (n_4013), .A (n_555));
XNOR2_X1 i_1416 (.ZN (n_4012), .A (n_4005), .B (n_4011));
XNOR2_X1 i_1415 (.ZN (n_4011), .A (n_282), .B (n_281));
AOI22_X1 i_1414 (.ZN (n_4005), .A1 (n_3934), .A2 (n_3935), .B1 (n_3933), .B2 (n_3932));
AOI22_X1 i_1413 (.ZN (n_4004), .A1 (n_3923), .A2 (n_4003), .B1 (n_4002), .B2 (n_4001));
XNOR2_X1 i_4050 (.ZN (result[46]), .A (n_3923), .B (n_4003));
XOR2_X1 i_1412 (.Z (n_4003), .A (n_4001), .B (n_4002));
AOI22_X1 i_1411 (.ZN (n_4002), .A1 (n_3919), .A2 (n_3884), .B1 (n_3886), .B2 (n_3918));
XNOR2_X1 i_1410 (.ZN (n_4001), .A (n_3957), .B (n_4000));
XOR2_X1 i_1409 (.Z (n_4000), .A (n_3997), .B (n_3999));
AOI22_X1 i_1408 (.ZN (n_3999), .A1 (n_3902), .A2 (n_3917), .B1 (n_3998), .B2 (n_3901));
INV_X1 i_1407 (.ZN (n_3998), .A (n_3887));
XOR2_X1 i_1406 (.Z (n_3997), .A (n_3995), .B (n_3996));
AOI22_X1 i_1405 (.ZN (n_3996), .A1 (n_3865), .A2 (n_3881), .B1 (n_3866), .B2 (n_3880));
XOR2_X1 i_1404 (.Z (n_3995), .A (n_3976), .B (n_3994));
XNOR2_X1 i_1403 (.ZN (n_3994), .A (n_546), .B (n_544));
OAI21_X1 i_1402 (.ZN (n_3976), .A (n_3975), .B1 (n_3958), .B2 (n_3974));
NAND2_X1 i_1401 (.ZN (n_3975), .A1 (n_3958), .A2 (n_3974));
XOR2_X1 i_1400 (.Z (n_3974), .A (n_3968), .B (n_551));
NAND2_X1 i_1399 (.ZN (n_3968), .A1 (n_561), .A2 (n_559));
AOI22_X1 i_1398 (.ZN (n_3958), .A1 (n_3899), .A2 (n_3900), .B1 (n_3893), .B2 (n_3898));
XOR2_X1 i_1397 (.Z (n_3957), .A (n_3954), .B (n_3956));
AOI22_X1 i_1396 (.ZN (n_3956), .A1 (n_3955), .A2 (n_3883), .B1 (n_3882), .B2 (n_3850));
INV_X1 i_1395 (.ZN (n_3955), .A (n_3849));
XOR2_X1 i_1394 (.Z (n_3954), .A (n_3931), .B (n_3953));
XNOR2_X1 i_1393 (.ZN (n_3953), .A (n_3943), .B (n_3952));
XNOR2_X1 i_1392 (.ZN (n_3952), .A (n_490), .B (n_486));
XOR2_X1 i_1391 (.Z (n_3943), .A (n_3936), .B (n_3942));
OAI21_X1 i_1390 (.ZN (n_3942), .A (n_442), .B1 (n_443), .B2 (n_445));
XNOR2_X1 i_1389 (.ZN (n_3936), .A (n_3934), .B (n_3935));
OAI21_X1 i_1388 (.ZN (n_3935), .A (n_3867), .B1 (n_3869), .B2 (n_509));
XOR2_X1 i_1387 (.Z (n_3934), .A (n_3932), .B (n_3933));
OAI33_X1 i_1386 (.ZN (n_3933), .A1 (n_3872), .A2 (n_217), .A3 (n_213), .B1 (n_389)
    , .B2 (n_216), .B3 (n_585));
OAI22_X1 i_1385 (.ZN (n_3932), .A1 (n_3877), .A2 (n_3878), .B1 (n_583), .B2 (n_3876));
XOR2_X1 i_1384 (.Z (n_3931), .A (n_3925), .B (n_3930));
XOR2_X1 i_1383 (.Z (n_3930), .A (n_3928), .B (n_3929));
AOI22_X1 i_1382 (.ZN (n_3929), .A1 (n_3851), .A2 (n_3864), .B1 (n_3857), .B2 (n_3863));
XNOR2_X1 i_1381 (.ZN (n_3928), .A (n_3926), .B (n_3927));
OAI22_X1 i_1380 (.ZN (n_3927), .A1 (n_3875), .A2 (n_3879), .B1 (n_3874), .B2 (n_3870));
AOI22_X1 i_1379 (.ZN (n_3926), .A1 (n_3905), .A2 (n_3910), .B1 (n_3904), .B2 (n_3903));
AOI22_X1 i_1378 (.ZN (n_3925), .A1 (n_3914), .A2 (n_3924), .B1 (n_3911), .B2 (n_3913));
INV_X1 i_1377 (.ZN (n_3924), .A (n_3916));
OAI22_X1 i_1376 (.ZN (n_3923), .A1 (n_3847), .A2 (n_3921), .B1 (n_3922), .B2 (n_3920));
INV_X1 i_1375 (.ZN (n_3922), .A (n_3848));
XNOR2_X1 i_3967 (.ZN (result[45]), .A (n_3847), .B (n_3921));
XOR2_X1 i_1374 (.Z (n_3921), .A (n_3848), .B (n_3920));
XOR2_X1 i_1373 (.Z (n_3920), .A (n_3884), .B (n_3919));
XOR2_X1 i_1372 (.Z (n_3919), .A (n_3886), .B (n_3918));
XNOR2_X1 i_1371 (.ZN (n_3918), .A (n_3902), .B (n_3917));
XNOR2_X1 i_1370 (.ZN (n_3917), .A (n_3914), .B (n_3916));
AOI22_X1 i_1369 (.ZN (n_3916), .A1 (n_3832), .A2 (n_3831), .B1 (n_3915), .B2 (n_3830));
INV_X1 i_1368 (.ZN (n_3915), .A (n_3829));
XOR2_X1 i_1367 (.Z (n_3914), .A (n_3911), .B (n_3913));
AOI22_X1 i_1366 (.ZN (n_3913), .A1 (n_3912), .A2 (n_3825), .B1 (n_3819), .B2 (n_3824));
INV_X1 i_1365 (.ZN (n_3912), .A (n_3815));
XNOR2_X1 i_1364 (.ZN (n_3911), .A (n_3905), .B (n_3910));
XOR2_X1 i_1363 (.Z (n_3910), .A (n_556), .B (n_574));
XOR2_X1 i_1362 (.Z (n_3905), .A (n_3903), .B (n_3904));
OAI21_X1 i_1361 (.ZN (n_3904), .A (n_3766), .B1 (n_3762), .B2 (n_3763));
OAI22_X1 i_1360 (.ZN (n_3903), .A1 (n_3772), .A2 (n_3773), .B1 (n_3769), .B2 (n_3771));
XNOR2_X1 i_1359 (.ZN (n_3902), .A (n_3887), .B (n_3901));
XNOR2_X1 i_1358 (.ZN (n_3901), .A (n_3899), .B (n_3900));
AOI22_X1 i_1357 (.ZN (n_3900), .A1 (n_3805), .A2 (n_3792), .B1 (n_3798), .B2 (n_3804));
XOR2_X1 i_1356 (.Z (n_3899), .A (n_3893), .B (n_3898));
XOR2_X1 i_1355 (.Z (n_3898), .A (n_495), .B (n_491));
XOR2_X1 i_1354 (.Z (n_3893), .A (n_571), .B (n_565));
AOI22_X1 i_1353 (.ZN (n_3887), .A1 (n_3808), .A2 (n_3807), .B1 (n_3564), .B2 (n_3806));
AOI22_X1 i_1352 (.ZN (n_3886), .A1 (n_3885), .A2 (n_3835), .B1 (n_3812), .B2 (n_3834));
INV_X1 i_1351 (.ZN (n_3885), .A (n_3837));
XOR2_X1 i_1350 (.Z (n_3884), .A (n_3849), .B (n_3883));
XOR2_X1 i_1349 (.Z (n_3883), .A (n_3850), .B (n_3882));
XNOR2_X1 i_1348 (.ZN (n_3882), .A (n_3865), .B (n_3881));
XOR2_X1 i_1347 (.Z (n_3881), .A (n_3866), .B (n_3880));
XNOR2_X1 i_1346 (.ZN (n_3880), .A (n_3875), .B (n_3879));
XOR2_X1 i_1345 (.Z (n_3879), .A (n_3877), .B (n_3878));
NAND2_X1 i_1344 (.ZN (n_3878), .A1 (inputB[19]), .A2 (inputA[26]));
XNOR2_X1 i_1343 (.ZN (n_3877), .A (n_583), .B (n_3876));
NAND2_X1 i_1342 (.ZN (n_3876), .A1 (inputB[17]), .A2 (inputA[28]));
XNOR2_X1 i_1341 (.ZN (n_3875), .A (n_3870), .B (n_3874));
XOR2_X1 i_1340 (.Z (n_3874), .A (n_3872), .B (n_3873));
NAND2_X1 i_1339 (.ZN (n_3873), .A1 (inputB[22]), .A2 (inputA[23]));
XNOR2_X1 i_1338 (.ZN (n_3872), .A (n_570), .B (n_389));
XOR2_X1 i_1337 (.Z (n_3870), .A (n_3869), .B (n_509));
NAND2_X1 i_1336 (.ZN (n_3869), .A1 (n_3867), .A2 (n_3868));
OAI22_X1 i_1335 (.ZN (n_3868), .A1 (n_482), .A2 (n_461), .B1 (n_259), .B2 (n_218));
NAND3_X1 i_1334 (.ZN (n_3867), .A1 (n_500), .A2 (inputA[22]), .A3 (inputB[24]));
AOI22_X1 i_1333 (.ZN (n_3866), .A1 (n_3779), .A2 (n_3767), .B1 (n_3774), .B2 (n_3778));
XOR2_X1 i_1332 (.Z (n_3865), .A (n_3851), .B (n_3864));
XOR2_X1 i_1331 (.Z (n_3864), .A (n_3857), .B (n_3863));
XOR2_X1 i_1330 (.Z (n_3863), .A (n_522), .B (n_521));
XOR2_X1 i_1329 (.Z (n_3857), .A (n_515), .B (n_514));
AOI22_X1 i_1328 (.ZN (n_3851), .A1 (n_3604), .A2 (n_3565), .B1 (n_3571), .B2 (n_3566));
OAI21_X1 i_1327 (.ZN (n_3850), .A (n_3827), .B1 (n_3828), .B2 (n_3833));
AOI22_X1 i_1326 (.ZN (n_3849), .A1 (n_3809), .A2 (n_3781), .B1 (n_3760), .B2 (n_3780));
AOI22_X1 i_1325 (.ZN (n_3848), .A1 (n_3811), .A2 (n_3838), .B1 (n_3759), .B2 (n_3810));
OAI21_X1 i_1324 (.ZN (n_3847), .A (n_3844), .B1 (n_3757), .B2 (n_3846));
NOR2_X1 i_1323 (.ZN (n_3846), .A1 (n_3839), .A2 (n_3845));
INV_X1 i_1322 (.ZN (n_3845), .A (n_3755));
OAI21_X1 i_1321 (.ZN (n_3844), .A (n_3840), .B1 (n_3660), .B2 (n_3843));
INV_X1 i_1320 (.ZN (n_3843), .A (n_3841));
XNOR2_X1 i_3887 (.ZN (result[44]), .A (n_3758), .B (n_3842));
NAND2_X1 i_3886 (.ZN (n_3842), .A1 (n_3840), .A2 (n_3841));
NAND2_X1 i_1319 (.ZN (n_3841), .A1 (n_3839), .A2 (n_3754));
OR2_X1 i_1318 (.ZN (n_3840), .A1 (n_3839), .A2 (n_3754));
XOR2_X1 i_1317 (.Z (n_3839), .A (n_3811), .B (n_3838));
XOR2_X1 i_1316 (.Z (n_3838), .A (n_3835), .B (n_3837));
AOI22_X1 i_1315 (.ZN (n_3837), .A1 (n_3728), .A2 (n_3752), .B1 (n_3836), .B2 (n_3727));
INV_X1 i_1314 (.ZN (n_3836), .A (n_3713));
XOR2_X1 i_1313 (.Z (n_3835), .A (n_3812), .B (n_3834));
XOR2_X1 i_1312 (.Z (n_3834), .A (n_3828), .B (n_3833));
XNOR2_X1 i_1311 (.ZN (n_3833), .A (n_3831), .B (n_3832));
AOI22_X1 i_1310 (.ZN (n_3832), .A1 (n_3799), .A2 (n_3791), .B1 (n_3871), .B2 (n_3800));
XNOR2_X1 i_1309 (.ZN (n_3831), .A (n_3829), .B (n_3830));
OAI21_X1 i_1308 (.ZN (n_3830), .A (n_3743), .B1 (n_3744), .B2 (n_3750));
AOI22_X1 i_1307 (.ZN (n_3829), .A1 (n_3695), .A2 (n_3702), .B1 (n_3688), .B2 (n_3694));
OAI21_X1 i_1306 (.ZN (n_3828), .A (n_3827), .B1 (n_3813), .B2 (n_3826));
NAND2_X1 i_1305 (.ZN (n_3827), .A1 (n_3813), .A2 (n_3826));
XOR2_X1 i_1304 (.Z (n_3826), .A (n_3815), .B (n_3825));
XOR2_X1 i_1303 (.Z (n_3825), .A (n_3819), .B (n_3824));
XOR2_X1 i_1302 (.Z (n_3824), .A (n_579), .B (n_578));
XOR2_X1 i_1301 (.Z (n_3819), .A (n_575), .B (n_3818));
NAND2_X1 i_1300 (.ZN (n_3818), .A1 (inputB[16]), .A2 (inputA[28]));
AOI22_X1 i_1299 (.ZN (n_3815), .A1 (n_3794), .A2 (n_3793), .B1 (n_3797), .B2 (n_3795));
AOI22_X1 i_1297 (.ZN (n_3813), .A1 (n_3790), .A2 (n_3888), .B1 (n_3896), .B2 (n_3889));
OAI22_X1 i_1296 (.ZN (n_3812), .A1 (n_3706), .A2 (n_3704), .B1 (n_3789), .B2 (n_3703));
XOR2_X1 i_1295 (.Z (n_3811), .A (n_3759), .B (n_3810));
XNOR2_X1 i_1294 (.ZN (n_3810), .A (n_3781), .B (n_3809));
XOR2_X1 i_1293 (.Z (n_3809), .A (n_3807), .B (n_3808));
AOI22_X1 i_1292 (.ZN (n_3808), .A1 (n_3720), .A2 (n_3726), .B1 (n_3714), .B2 (n_3719));
XOR2_X1 i_1291 (.Z (n_3807), .A (n_3564), .B (n_3806));
XOR2_X1 i_1290 (.Z (n_3806), .A (n_3792), .B (n_3805));
XOR2_X1 i_1289 (.Z (n_3805), .A (n_3798), .B (n_3804));
XNOR2_X1 i_1288 (.ZN (n_3804), .A (n_506), .B (n_500));
XNOR2_X1 i_1287 (.ZN (n_3798), .A (n_567), .B (n_566));
XNOR2_X1 i_1286 (.ZN (n_3792), .A (n_512), .B (n_511));
XOR2_X1 i_1285 (.Z (n_3781), .A (n_3760), .B (n_3780));
XOR2_X1 i_1284 (.Z (n_3780), .A (n_3767), .B (n_3779));
XOR2_X1 i_1283 (.Z (n_3779), .A (n_3774), .B (n_3778));
XNOR2_X1 i_1282 (.ZN (n_3778), .A (n_493), .B (n_492));
XNOR2_X1 i_1281 (.ZN (n_3774), .A (n_3772), .B (n_3773));
AOI21_X1 i_1280 (.ZN (n_3773), .A (n_3746), .B1 (n_3748), .B2 (n_3749));
AOI22_X1 i_1279 (.ZN (n_3772), .A1 (n_3769), .A2 (n_3770), .B1 (n_3771), .B2 (n_3768));
INV_X1 i_1278 (.ZN (n_3771), .A (n_3770));
OAI21_X1 i_1277 (.ZN (n_3770), .A (n_3699), .B1 (n_3700), .B2 (n_3701));
INV_X1 i_1276 (.ZN (n_3769), .A (n_3768));
OAI22_X1 i_1275 (.ZN (n_3768), .A1 (n_3741), .A2 (n_3596), .B1 (n_510), .B2 (n_3740));
OAI21_X1 i_1274 (.ZN (n_3767), .A (n_3766), .B1 (n_3765), .B2 (n_3764));
NAND2_X1 i_1273 (.ZN (n_3766), .A1 (n_3764), .A2 (n_3765));
NAND2_X1 i_1272 (.ZN (n_3765), .A1 (inputB[13]), .A2 (inputA[31]));
XOR2_X1 i_1271 (.Z (n_3764), .A (n_3762), .B (n_3763));
AOI21_X1 i_1270 (.ZN (n_3763), .A (n_3690), .B1 (n_3692), .B2 (n_3693));
AOI21_X1 i_1269 (.ZN (n_3762), .A (n_3684), .B1 (n_3686), .B2 (n_3761));
INV_X1 i_1268 (.ZN (n_3761), .A (n_584));
AOI22_X1 i_1267 (.ZN (n_3760), .A1 (n_3732), .A2 (n_3751), .B1 (n_3626), .B2 (n_3730));
AOI22_X1 i_1266 (.ZN (n_3759), .A1 (n_3667), .A2 (n_3708), .B1 (n_3668), .B2 (n_3707));
NAND2_X1 i_3802 (.ZN (n_3758), .A1 (n_3661), .A2 (n_3757));
NAND2_X1 i_1265 (.ZN (n_3757), .A1 (n_3662), .A2 (n_3756));
XNOR2_X1 i_3800 (.ZN (result[43]), .A (n_3663), .B (n_3756));
AOI22_X1 i_1264 (.ZN (n_3756), .A1 (n_3754), .A2 (n_3755), .B1 (n_3711), .B2 (n_3753));
OR2_X1 i_1263 (.ZN (n_3755), .A1 (n_3710), .A2 (n_3753));
OAI21_X1 i_1262 (.ZN (n_3754), .A (n_3710), .B1 (n_3711), .B2 (n_3753));
XOR2_X1 i_1261 (.Z (n_3753), .A (n_3728), .B (n_3752));
XNOR2_X1 i_1260 (.ZN (n_3752), .A (n_3732), .B (n_3751));
XNOR2_X1 i_1259 (.ZN (n_3751), .A (n_3744), .B (n_3750));
XOR2_X1 i_1258 (.Z (n_3750), .A (n_3748), .B (n_3749));
NOR2_X1 i_1257 (.ZN (n_3749), .A1 (n_478), .A2 (n_127));
NOR2_X1 i_1256 (.ZN (n_3748), .A1 (n_3746), .A2 (n_3747));
AOI22_X1 i_1255 (.ZN (n_3747), .A1 (inputA[17]), .A2 (inputB[26]), .B1 (inputA[16]), .B2 (inputB[27]));
NOR2_X1 i_1254 (.ZN (n_3746), .A1 (n_3602), .A2 (n_513));
OAI21_X1 i_1253 (.ZN (n_3744), .A (n_3743), .B1 (n_3738), .B2 (n_3742));
NAND2_X1 i_1252 (.ZN (n_3743), .A1 (n_3738), .A2 (n_3742));
XNOR2_X1 i_1251 (.ZN (n_3742), .A (n_3741), .B (n_3596));
XNOR2_X1 i_1250 (.ZN (n_3741), .A (n_510), .B (n_3740));
NAND2_X1 i_1249 (.ZN (n_3740), .A1 (inputA[20]), .A2 (inputB[23]));
XNOR2_X1 i_1248 (.ZN (n_3738), .A (n_3568), .B (n_3567));
XOR2_X1 i_1247 (.Z (n_3732), .A (n_3730), .B (n_3626));
AOI22_X1 i_1246 (.ZN (n_3730), .A1 (n_3644), .A2 (n_3729), .B1 (n_3635), .B2 (n_3643));
INV_X1 i_1245 (.ZN (n_3729), .A (n_3645));
XNOR2_X1 i_1244 (.ZN (n_3728), .A (n_3713), .B (n_3727));
XNOR2_X1 i_1243 (.ZN (n_3727), .A (n_3720), .B (n_3726));
XOR2_X1 i_1242 (.Z (n_3726), .A (n_3610), .B (n_3605));
XOR2_X1 i_1241 (.Z (n_3720), .A (n_3714), .B (n_3719));
XOR2_X1 i_1240 (.Z (n_3719), .A (n_3588), .B (n_3572));
OAI22_X1 i_1239 (.ZN (n_3714), .A1 (n_4244), .A2 (n_4220), .B1 (n_4227), .B2 (n_4221));
AOI22_X1 i_1238 (.ZN (n_3713), .A1 (n_3600), .A2 (n_3614), .B1 (n_3712), .B2 (n_3599));
INV_X1 i_1237 (.ZN (n_3712), .A (n_3583));
NOR2_X1 i_1236 (.ZN (n_3711), .A1 (n_3665), .A2 (n_3709));
NAND2_X1 i_1235 (.ZN (n_3710), .A1 (n_3665), .A2 (n_3709));
XNOR2_X1 i_1234 (.ZN (n_3709), .A (n_3667), .B (n_3708));
XOR2_X1 i_1233 (.Z (n_3708), .A (n_3668), .B (n_3707));
XOR2_X1 i_1232 (.Z (n_3707), .A (n_3704), .B (n_3706));
AOI22_X1 i_1231 (.ZN (n_3706), .A1 (n_4164), .A2 (n_3705), .B1 (n_4218), .B2 (n_4165));
INV_X1 i_1230 (.ZN (n_3705), .A (n_3574));
XNOR2_X1 i_1229 (.ZN (n_3704), .A (n_3789), .B (n_3703));
XNOR2_X1 i_1228 (.ZN (n_3703), .A (n_3695), .B (n_3702));
XNOR2_X1 i_1227 (.ZN (n_3702), .A (n_3700), .B (n_3701));
NAND2_X1 i_1226 (.ZN (n_3701), .A1 (inputA[21]), .A2 (inputB[22]));
OAI21_X1 i_1225 (.ZN (n_3700), .A (n_3699), .B1 (n_3696), .B2 (n_3698));
NAND2_X1 i_1224 (.ZN (n_3699), .A1 (n_3696), .A2 (n_3698));
NOR2_X1 i_1223 (.ZN (n_3698), .A1 (n_216), .A2 (n_259));
NOR2_X1 i_1222 (.ZN (n_3696), .A1 (n_414), .A2 (n_213));
XOR2_X1 i_1221 (.Z (n_3695), .A (n_3688), .B (n_3694));
XNOR2_X1 i_1220 (.ZN (n_3694), .A (n_3692), .B (n_3693));
NOR2_X1 i_1219 (.ZN (n_3693), .A1 (n_588), .A2 (n_215));
NOR2_X1 i_1218 (.ZN (n_3692), .A1 (n_3690), .A2 (n_3691));
AOI22_X1 i_1217 (.ZN (n_3691), .A1 (inputB[14]), .A2 (inputA[29]), .B1 (inputB[15]), .B2 (inputA[28]));
NOR2_X1 i_1216 (.ZN (n_3690), .A1 (n_3624), .A2 (n_577));
XOR2_X1 i_1215 (.Z (n_3688), .A (n_3686), .B (n_584));
NOR2_X1 i_1214 (.ZN (n_3686), .A1 (n_3684), .A2 (n_3685));
AOI22_X1 i_1213 (.ZN (n_3685), .A1 (inputB[18]), .A2 (inputA[25]), .B1 (inputB[19]), .B2 (inputA[24]));
NOR3_X1 i_1212 (.ZN (n_3684), .A1 (n_578), .A2 (n_400), .A3 (n_585));
AOI22_X1 i_1211 (.ZN (n_3668), .A1 (n_3634), .A2 (n_3646), .B1 (n_3617), .B2 (n_3633));
AOI22_X1 i_1210 (.ZN (n_3667), .A1 (n_3576), .A2 (n_3578), .B1 (n_3666), .B2 (n_3575));
INV_X1 i_1209 (.ZN (n_3666), .A (n_4275));
OAI22_X1 i_1208 (.ZN (n_3665), .A1 (n_3664), .A2 (n_3648), .B1 (n_3647), .B2 (n_3615));
INV_X1 i_1207 (.ZN (n_3664), .A (n_3581));
NAND2_X1 i_3706 (.ZN (n_3663), .A1 (n_3661), .A2 (n_3662));
NAND2_X1 i_1206 (.ZN (n_3662), .A1 (n_3656), .A2 (n_3659));
INV_X1 i_3704 (.ZN (n_3661), .A (n_3660));
NOR2_X1 i_1205 (.ZN (n_3660), .A1 (n_3656), .A2 (n_3659));
AOI21_X1 i_1204 (.ZN (n_3659), .A (n_3657), .B1 (n_3658), .B2 (n_3579));
INV_X1 i_1203 (.ZN (n_3658), .A (n_3561));
INV_X1 i_1202 (.ZN (n_3657), .A (n_3650));
OAI22_X1 i_1201 (.ZN (n_3656), .A1 (n_3559), .A2 (n_3654), .B1 (n_3655), .B2 (n_3653));
INV_X1 i_1200 (.ZN (n_3655), .A (n_3651));
XNOR2_X1 i_3697 (.ZN (result[42]), .A (n_3559), .B (n_3654));
XOR2_X1 i_1199 (.Z (n_3654), .A (n_3651), .B (n_3653));
AOI22_X1 i_1198 (.ZN (n_3653), .A1 (n_3527), .A2 (n_3555), .B1 (n_3652), .B2 (n_3554));
INV_X1 i_1197 (.ZN (n_3652), .A (n_3529));
OAI21_X1 i_1196 (.ZN (n_3651), .A (n_3650), .B1 (n_3580), .B2 (n_3649));
NAND2_X1 i_1195 (.ZN (n_3650), .A1 (n_3580), .A2 (n_3649));
XNOR2_X1 i_1194 (.ZN (n_3649), .A (n_3581), .B (n_3648));
XNOR2_X1 i_1193 (.ZN (n_3648), .A (n_3615), .B (n_3647));
XNOR2_X1 i_1192 (.ZN (n_3647), .A (n_3634), .B (n_3646));
XOR2_X1 i_1191 (.Z (n_3646), .A (n_3644), .B (n_3645));
AOI22_X1 i_1190 (.ZN (n_3645), .A1 (n_4287), .A2 (n_4286), .B1 (n_4289), .B2 (n_4288));
XOR2_X1 i_1189 (.Z (n_3644), .A (n_3635), .B (n_3643));
XNOR2_X1 i_1188 (.ZN (n_3643), .A (n_3821), .B (n_3801));
AOI22_X1 i_1187 (.ZN (n_3635), .A1 (n_4279), .A2 (n_4285), .B1 (n_4280), .B2 (n_4282));
XOR2_X1 i_1186 (.Z (n_3634), .A (n_3617), .B (n_3633));
XNOR2_X1 i_1185 (.ZN (n_3633), .A (n_3721), .B (n_3627));
AOI22_X1 i_1184 (.ZN (n_3617), .A1 (n_3549), .A2 (n_3616), .B1 (n_3548), .B2 (n_3546));
INV_X1 i_1183 (.ZN (n_3616), .A (n_3551));
XOR2_X1 i_1182 (.Z (n_3615), .A (n_3600), .B (n_3614));
XOR2_X1 i_1181 (.Z (n_3614), .A (n_3907), .B (n_3897));
XNOR2_X1 i_1180 (.ZN (n_3600), .A (n_3583), .B (n_3599));
XOR2_X1 i_1179 (.Z (n_3599), .A (n_3891), .B (n_3890));
AOI22_X1 i_1178 (.ZN (n_3583), .A1 (n_3505), .A2 (n_3513), .B1 (n_3502), .B2 (n_3582));
INV_X1 i_1177 (.ZN (n_3582), .A (n_3504));
AOI22_X1 i_1176 (.ZN (n_3581), .A1 (n_3531), .A2 (n_3553), .B1 (n_3533), .B2 (n_3552));
XNOR2_X1 i_1175 (.ZN (n_3580), .A (n_3561), .B (n_3579));
XOR2_X1 i_1174 (.Z (n_3579), .A (n_3576), .B (n_3578));
AOI22_X1 i_1173 (.ZN (n_3578), .A1 (n_3577), .A2 (n_3524), .B1 (n_3514), .B2 (n_3523));
INV_X1 i_1172 (.ZN (n_3577), .A (n_3944));
XNOR2_X1 i_1171 (.ZN (n_3576), .A (n_4275), .B (n_3575));
XOR2_X1 i_1170 (.Z (n_3575), .A (n_4164), .B (n_3574));
AOI22_X1 i_1169 (.ZN (n_3574), .A1 (n_3573), .A2 (n_3522), .B1 (n_3521), .B2 (n_3520));
INV_X1 i_1168 (.ZN (n_3573), .A (n_3515));
AOI22_X1 i_1167 (.ZN (n_3561), .A1 (n_3495), .A2 (n_3526), .B1 (n_3560), .B2 (n_3494));
INV_X1 i_1166 (.ZN (n_3560), .A (n_3450));
AOI22_X1 i_1165 (.ZN (n_3559), .A1 (n_3447), .A2 (n_3558), .B1 (n_3556), .B2 (n_3557));
XNOR2_X1 i_3600 (.ZN (result[41]), .A (n_3447), .B (n_3558));
XOR2_X1 i_1164 (.Z (n_3558), .A (n_3556), .B (n_3557));
OAI21_X1 i_1163 (.ZN (n_3557), .A (n_3443), .B1 (n_3366), .B2 (n_3365));
XOR2_X1 i_1162 (.Z (n_3556), .A (n_3527), .B (n_3555));
XNOR2_X1 i_1161 (.ZN (n_3555), .A (n_3529), .B (n_3554));
XOR2_X1 i_1160 (.Z (n_3554), .A (n_3531), .B (n_3553));
XOR2_X1 i_1159 (.Z (n_3553), .A (n_3533), .B (n_3552));
XNOR2_X1 i_1158 (.ZN (n_3552), .A (n_3549), .B (n_3551));
AOI22_X1 i_1157 (.ZN (n_3551), .A1 (n_3435), .A2 (n_3550), .B1 (n_3434), .B2 (n_3427));
INV_X1 i_1156 (.ZN (n_3550), .A (n_3436));
XOR2_X1 i_1155 (.Z (n_3549), .A (n_3546), .B (n_3548));
AOI22_X1 i_1154 (.ZN (n_3548), .A1 (n_3547), .A2 (n_3949), .B1 (n_3950), .B2 (n_3951));
INV_X1 i_1153 (.ZN (n_3547), .A (n_3948));
XNOR2_X1 i_1152 (.ZN (n_3546), .A (n_4192), .B (n_4168));
AOI22_X1 i_1151 (.ZN (n_3533), .A1 (n_3532), .A2 (n_3404), .B1 (n_3385), .B2 (n_3403));
INV_X1 i_1150 (.ZN (n_3532), .A (n_3369));
AOI22_X1 i_1149 (.ZN (n_3531), .A1 (n_3438), .A2 (n_3530), .B1 (n_3419), .B2 (n_3437));
INV_X1 i_1148 (.ZN (n_3530), .A (n_3406));
AOI22_X1 i_1147 (.ZN (n_3529), .A1 (n_3440), .A2 (n_3528), .B1 (n_3439), .B2 (n_3405));
INV_X1 i_1146 (.ZN (n_3528), .A (n_3441));
XNOR2_X1 i_1145 (.ZN (n_3527), .A (n_3495), .B (n_3526));
XOR2_X1 i_1144 (.Z (n_3526), .A (n_3524), .B (n_3944));
XOR2_X1 i_1143 (.Z (n_3524), .A (n_3514), .B (n_3523));
XNOR2_X1 i_1142 (.ZN (n_3523), .A (n_3515), .B (n_3522));
XOR2_X1 i_1141 (.Z (n_3522), .A (n_3520), .B (n_3521));
OAI21_X1 i_1140 (.ZN (n_3521), .A (n_3402), .B1 (n_3395), .B2 (n_3389));
XNOR2_X1 i_1139 (.ZN (n_3520), .A (n_4238), .B (n_4232));
AOI22_X1 i_1138 (.ZN (n_3515), .A1 (n_3380), .A2 (n_3384), .B1 (n_3375), .B2 (n_3379));
XOR2_X1 i_1137 (.Z (n_3514), .A (n_3505), .B (n_3513));
XOR2_X1 i_1136 (.Z (n_3513), .A (n_3642), .B (n_3628));
XNOR2_X1 i_1135 (.ZN (n_3505), .A (n_3502), .B (n_3504));
AOI22_X1 i_1134 (.ZN (n_3504), .A1 (n_4293), .A2 (n_4292), .B1 (n_3503), .B2 (n_4294));
INV_X1 i_1133 (.ZN (n_3503), .A (n_4295));
XOR2_X1 i_1132 (.Z (n_3502), .A (n_4256), .B (n_4245));
XNOR2_X1 i_1131 (.ZN (n_3495), .A (n_3450), .B (n_3494));
XOR2_X1 i_1130 (.Z (n_3494), .A (n_4290), .B (n_4276));
AOI22_X1 i_1129 (.ZN (n_3450), .A1 (n_3363), .A2 (n_3448), .B1 (n_3449), .B2 (n_3362));
INV_X1 i_1128 (.ZN (n_3449), .A (n_3345));
INV_X1 i_1127 (.ZN (n_3448), .A (n_3364));
OAI22_X1 i_1126 (.ZN (n_3447), .A1 (n_3343), .A2 (n_3445), .B1 (n_3446), .B2 (n_3444));
INV_X1 i_1125 (.ZN (n_3446), .A (n_3344));
XNOR2_X1 i_3486 (.ZN (result[40]), .A (n_3343), .B (n_3445));
XOR2_X1 i_1124 (.Z (n_3445), .A (n_3344), .B (n_3444));
OAI21_X1 i_1123 (.ZN (n_3444), .A (n_3443), .B1 (n_3367), .B2 (n_3442));
NAND2_X1 i_1122 (.ZN (n_3443), .A1 (n_3367), .A2 (n_3442));
XNOR2_X1 i_1121 (.ZN (n_3442), .A (n_3440), .B (n_3441));
AOI22_X1 i_1120 (.ZN (n_3441), .A1 (n_3333), .A2 (n_3307), .B1 (n_3308), .B2 (n_3332));
XOR2_X1 i_1119 (.Z (n_3440), .A (n_3405), .B (n_3439));
XOR2_X1 i_1118 (.Z (n_3439), .A (n_3406), .B (n_3438));
XOR2_X1 i_1117 (.Z (n_3438), .A (n_3419), .B (n_3437));
XOR2_X1 i_1116 (.Z (n_3437), .A (n_3435), .B (n_3436));
AOI22_X1 i_1115 (.ZN (n_3436), .A1 (n_3322), .A2 (n_3328), .B1 (n_3317), .B2 (n_3321));
XOR2_X1 i_1114 (.Z (n_3435), .A (n_3427), .B (n_3434));
XNOR2_X1 i_1113 (.ZN (n_3434), .A (n_4175), .B (n_4169));
XOR2_X1 i_1112 (.Z (n_3427), .A (n_3677), .B (n_3670));
XNOR2_X1 i_1111 (.ZN (n_3419), .A (n_4296), .B (n_4291));
AOI22_X1 i_1110 (.ZN (n_3406), .A1 (n_3330), .A2 (n_3331), .B1 (n_3311), .B2 (n_3329));
XOR2_X1 i_1109 (.Z (n_3405), .A (n_3369), .B (n_3404));
XOR2_X1 i_1108 (.Z (n_3404), .A (n_3385), .B (n_3403));
OAI21_X1 i_1107 (.ZN (n_3403), .A (n_3402), .B1 (n_3401), .B2 (n_3396));
NAND2_X1 i_1106 (.ZN (n_3402), .A1 (n_3396), .A2 (n_3401));
XOR2_X1 i_1105 (.Z (n_3401), .A (n_4248), .B (n_3689));
XOR2_X1 i_1104 (.Z (n_3396), .A (n_3389), .B (n_3395));
XOR2_X1 i_1103 (.Z (n_3395), .A (n_4261), .B (n_3788));
XOR2_X1 i_1102 (.Z (n_3389), .A (n_4259), .B (n_3388));
NAND2_X1 i_1101 (.ZN (n_3388), .A1 (inputB[19]), .A2 (inputA[21]));
XNOR2_X1 i_1100 (.ZN (n_3385), .A (n_3380), .B (n_3384));
XNOR2_X1 i_1099 (.ZN (n_3384), .A (n_4242), .B (n_4241));
XOR2_X1 i_1098 (.Z (n_3380), .A (n_3375), .B (n_3379));
XNOR2_X1 i_1097 (.ZN (n_3379), .A (n_4234), .B (n_4233));
XNOR2_X1 i_1096 (.ZN (n_3375), .A (n_4197), .B (n_4196));
AOI22_X1 i_1095 (.ZN (n_3369), .A1 (n_3241), .A2 (n_3368), .B1 (n_3239), .B2 (n_3240));
INV_X1 i_1094 (.ZN (n_3368), .A (n_3242));
XOR2_X1 i_1093 (.Z (n_3367), .A (n_3365), .B (n_3366));
AOI22_X1 i_1092 (.ZN (n_3366), .A1 (n_3264), .A2 (n_3266), .B1 (n_3261), .B2 (n_3263));
XNOR2_X1 i_1091 (.ZN (n_3365), .A (n_3363), .B (n_3364));
AOI22_X1 i_1090 (.ZN (n_3364), .A1 (n_3305), .A2 (n_3306), .B1 (n_3282), .B2 (n_3304));
XNOR2_X1 i_1089 (.ZN (n_3363), .A (n_3345), .B (n_3362));
XNOR2_X1 i_1088 (.ZN (n_3362), .A (n_4034), .B (n_3945));
AOI22_X1 i_1087 (.ZN (n_3345), .A1 (n_3258), .A2 (n_3260), .B1 (n_3243), .B2 (n_3257));
OAI21_X1 i_1086 (.ZN (n_3344), .A (n_3338), .B1 (n_3267), .B2 (n_3334));
AOI22_X1 i_1085 (.ZN (n_3343), .A1 (n_3231), .A2 (n_3341), .B1 (n_3342), .B2 (n_3340));
INV_X1 i_1084 (.ZN (n_3342), .A (n_3339));
XNOR2_X1 i_3381 (.ZN (result[39]), .A (n_3231), .B (n_3341));
XNOR2_X1 i_1083 (.ZN (n_3341), .A (n_3339), .B (n_3340));
OAI22_X1 i_1082 (.ZN (n_3340), .A1 (n_3190), .A2 (n_3228), .B1 (n_3126), .B2 (n_3189));
OAI21_X1 i_1081 (.ZN (n_3339), .A (n_3338), .B1 (n_3335), .B2 (n_3337));
NAND2_X1 i_1080 (.ZN (n_3338), .A1 (n_3335), .A2 (n_3337));
AOI22_X1 i_1079 (.ZN (n_3337), .A1 (n_3336), .A2 (n_3226), .B1 (n_3191), .B2 (n_3225));
INV_X1 i_1078 (.ZN (n_3336), .A (n_3227));
XOR2_X1 i_1077 (.Z (n_3335), .A (n_3267), .B (n_3334));
XNOR2_X1 i_1076 (.ZN (n_3334), .A (n_3307), .B (n_3333));
XOR2_X1 i_1075 (.Z (n_3333), .A (n_3308), .B (n_3332));
XNOR2_X1 i_1074 (.ZN (n_3332), .A (n_3330), .B (n_3331));
AOI22_X1 i_1073 (.ZN (n_3331), .A1 (n_3203), .A2 (n_3210), .B1 (n_3197), .B2 (n_3202));
XOR2_X1 i_1072 (.Z (n_3330), .A (n_3311), .B (n_3329));
XNOR2_X1 i_1071 (.ZN (n_3329), .A (n_3322), .B (n_3328));
XNOR2_X1 i_1070 (.ZN (n_3328), .A (n_3672), .B (n_3671));
XOR2_X1 i_1069 (.Z (n_3322), .A (n_3317), .B (n_3321));
XNOR2_X1 i_1068 (.ZN (n_3321), .A (n_3716), .B (n_3715));
XOR2_X1 i_1067 (.Z (n_3317), .A (n_3681), .B (n_3680));
AOI22_X1 i_1066 (.ZN (n_3311), .A1 (n_3309), .A2 (n_3166), .B1 (n_3310), .B2 (n_3164));
INV_X1 i_1065 (.ZN (n_3310), .A (n_3165));
INV_X1 i_1064 (.ZN (n_3309), .A (n_3163));
OAI22_X1 i_1063 (.ZN (n_3308), .A1 (n_3161), .A2 (n_3187), .B1 (n_3167), .B2 (n_3186));
XNOR2_X1 i_1062 (.ZN (n_3307), .A (n_3305), .B (n_3306));
AOI22_X1 i_1061 (.ZN (n_3306), .A1 (n_3221), .A2 (n_3223), .B1 (n_3219), .B2 (n_3220));
XOR2_X1 i_1060 (.Z (n_3305), .A (n_3282), .B (n_3304));
OAI21_X1 i_1059 (.ZN (n_3304), .A (n_4301), .B1 (n_4303), .B2 (n_4302));
XOR2_X1 i_1058 (.Z (n_3282), .A (n_4086), .B (n_4035));
XNOR2_X1 i_1057 (.ZN (n_3267), .A (n_3264), .B (n_3266));
AOI22_X1 i_1056 (.ZN (n_3266), .A1 (n_3160), .A2 (n_3188), .B1 (n_3265), .B2 (n_3159));
INV_X1 i_1055 (.ZN (n_3265), .A (n_3128));
XOR2_X1 i_1054 (.Z (n_3264), .A (n_3261), .B (n_3263));
AOI22_X1 i_1053 (.ZN (n_3263), .A1 (n_3212), .A2 (n_3224), .B1 (n_3262), .B2 (n_3211));
INV_X1 i_1052 (.ZN (n_3262), .A (n_3192));
XNOR2_X1 i_1051 (.ZN (n_3261), .A (n_3258), .B (n_3260));
AOI22_X1 i_1050 (.ZN (n_3260), .A1 (n_3143), .A2 (n_3158), .B1 (n_3259), .B2 (n_3142));
INV_X1 i_1049 (.ZN (n_3259), .A (n_3129));
XOR2_X1 i_1048 (.Z (n_3258), .A (n_3243), .B (n_3257));
XOR2_X1 i_1047 (.Z (n_3257), .A (n_3965), .B (n_3959));
XNOR2_X1 i_1046 (.ZN (n_3243), .A (n_3241), .B (n_3242));
AOI22_X1 i_1045 (.ZN (n_3242), .A1 (n_3130), .A2 (n_3141), .B1 (n_3140), .B2 (n_3135));
XOR2_X1 i_1044 (.Z (n_3241), .A (n_3239), .B (n_3240));
AOI22_X1 i_1043 (.ZN (n_3240), .A1 (n_3181), .A2 (n_3185), .B1 (n_3173), .B2 (n_3180));
XNOR2_X1 i_1042 (.ZN (n_3239), .A (n_4312), .B (n_4311));
OAI22_X1 i_1041 (.ZN (n_3231), .A1 (n_3124), .A2 (n_3230), .B1 (n_3125), .B2 (n_3229));
XNOR2_X1 i_3269 (.ZN (result[38]), .A (n_3124), .B (n_3230));
XNOR2_X1 i_1040 (.ZN (n_3230), .A (n_3125), .B (n_3229));
XNOR2_X1 i_1039 (.ZN (n_3229), .A (n_3190), .B (n_3228));
XNOR2_X1 i_1038 (.ZN (n_3228), .A (n_3226), .B (n_3227));
AOI22_X1 i_1037 (.ZN (n_3227), .A1 (n_3055), .A2 (n_3056), .B1 (n_3005), .B2 (n_3054));
XOR2_X1 i_1036 (.Z (n_3226), .A (n_3191), .B (n_3225));
XOR2_X1 i_1035 (.Z (n_3225), .A (n_3212), .B (n_3224));
XNOR2_X1 i_1034 (.ZN (n_3224), .A (n_3221), .B (n_3223));
AOI22_X1 i_1033 (.ZN (n_3223), .A1 (n_3091), .A2 (n_3092), .B1 (n_3222), .B2 (n_3089));
INV_X1 i_1032 (.ZN (n_3222), .A (n_3090));
XOR2_X1 i_1031 (.Z (n_3221), .A (n_3219), .B (n_3220));
AOI22_X1 i_1030 (.ZN (n_3220), .A1 (n_3006), .A2 (n_3015), .B1 (n_3010), .B2 (n_3014));
XNOR2_X1 i_1029 (.ZN (n_3219), .A (n_4112), .B (n_4097));
XNOR2_X1 i_1028 (.ZN (n_3212), .A (n_3192), .B (n_3211));
XNOR2_X1 i_1027 (.ZN (n_3211), .A (n_3203), .B (n_3210));
XNOR2_X1 i_1026 (.ZN (n_3210), .A (n_4321), .B (n_4316));
XOR2_X1 i_1025 (.Z (n_3203), .A (n_3197), .B (n_3202));
XNOR2_X1 i_1024 (.ZN (n_3202), .A (n_4061), .B (n_4042));
XNOR2_X1 i_1023 (.ZN (n_3197), .A (n_4364), .B (n_4350));
AOI22_X1 i_1022 (.ZN (n_3192), .A1 (n_3037), .A2 (n_3053), .B1 (n_3016), .B2 (n_3036));
OAI21_X1 i_1021 (.ZN (n_3191), .A (n_3084), .B1 (n_3063), .B2 (n_3064));
XNOR2_X1 i_1020 (.ZN (n_3190), .A (n_3126), .B (n_3189));
XOR2_X1 i_1019 (.Z (n_3189), .A (n_3160), .B (n_3188));
XNOR2_X1 i_1018 (.ZN (n_3188), .A (n_3161), .B (n_3187));
XNOR2_X1 i_1017 (.ZN (n_3187), .A (n_3167), .B (n_3186));
XNOR2_X1 i_1016 (.ZN (n_3186), .A (n_3181), .B (n_3185));
XNOR2_X1 i_1015 (.ZN (n_3185), .A (n_3971), .B (n_3970));
XOR2_X1 i_1014 (.Z (n_3181), .A (n_3173), .B (n_3180));
XNOR2_X1 i_1013 (.ZN (n_3180), .A (n_3980), .B (n_3979));
XOR2_X1 i_1012 (.Z (n_3173), .A (n_3988), .B (n_3987));
XOR2_X1 i_1011 (.Z (n_3167), .A (n_3163), .B (n_3166));
XNOR2_X1 i_1010 (.ZN (n_3166), .A (n_3164), .B (n_3165));
AOI22_X1 i_1009 (.ZN (n_3165), .A1 (n_3046), .A2 (n_3052), .B1 (n_3041), .B2 (n_3045));
OAI21_X1 i_1008 (.ZN (n_3164), .A (n_3035), .B1 (n_3027), .B2 (n_3021));
AOI22_X1 i_1007 (.ZN (n_3163), .A1 (n_3070), .A2 (n_3076), .B1 (n_3068), .B2 (n_3162));
INV_X1 i_1006 (.ZN (n_3162), .A (n_3069));
OAI21_X1 i_1005 (.ZN (n_3161), .A (n_3081), .B1 (n_3067), .B2 (n_3082));
XNOR2_X1 i_1004 (.ZN (n_3160), .A (n_3128), .B (n_3159));
XNOR2_X1 i_1003 (.ZN (n_3159), .A (n_3143), .B (n_3158));
XOR2_X1 i_1002 (.Z (n_3158), .A (n_3961), .B (n_3960));
XNOR2_X1 i_1001 (.ZN (n_3143), .A (n_3129), .B (n_3142));
XNOR2_X1 i_1000 (.ZN (n_3142), .A (n_3130), .B (n_3141));
XOR2_X1 i_999 (.Z (n_3141), .A (n_3135), .B (n_3140));
XOR2_X1 i_998 (.Z (n_3140), .A (n_4065), .B (n_3139));
NAND2_X1 i_997 (.ZN (n_3139), .A1 (inputA[10]), .A2 (inputB[28]));
XOR2_X1 i_996 (.Z (n_3135), .A (n_4082), .B (n_4067));
OAI22_X1 i_995 (.ZN (n_3130), .A1 (n_3112), .A2 (n_3115), .B1 (n_3113), .B2 (n_3114));
AOI22_X1 i_994 (.ZN (n_3129), .A1 (n_3109), .A2 (n_3116), .B1 (n_3100), .B2 (n_3108));
AOI22_X1 i_993 (.ZN (n_3128), .A1 (n_3094), .A2 (n_3117), .B1 (n_3127), .B2 (n_3093));
INV_X1 i_992 (.ZN (n_3127), .A (n_3088));
AOI22_X1 i_991 (.ZN (n_3126), .A1 (n_3119), .A2 (n_3062), .B1 (n_3085), .B2 (n_3118));
AOI22_X1 i_990 (.ZN (n_3125), .A1 (n_3060), .A2 (n_3120), .B1 (n_3059), .B2 (n_3057));
AOI22_X1 i_989 (.ZN (n_3124), .A1 (n_3004), .A2 (n_3123), .B1 (n_3121), .B2 (n_3122));
XNOR2_X1 i_3161 (.ZN (result[37]), .A (n_3004), .B (n_3123));
XOR2_X1 i_988 (.Z (n_3123), .A (n_3121), .B (n_3122));
OAI21_X1 i_987 (.ZN (n_3122), .A (n_2920), .B1 (n_2921), .B2 (n_3002));
XOR2_X1 i_986 (.Z (n_3121), .A (n_3060), .B (n_3120));
XOR2_X1 i_985 (.Z (n_3120), .A (n_3062), .B (n_3119));
XOR2_X1 i_984 (.Z (n_3119), .A (n_3085), .B (n_3118));
XNOR2_X1 i_983 (.ZN (n_3118), .A (n_3094), .B (n_3117));
XNOR2_X1 i_982 (.ZN (n_3117), .A (n_3109), .B (n_3116));
XNOR2_X1 i_981 (.ZN (n_3116), .A (n_3112), .B (n_3115));
XNOR2_X1 i_980 (.ZN (n_3115), .A (n_3113), .B (n_3114));
AOI21_X1 i_979 (.ZN (n_3114), .A (n_2991), .B1 (n_2993), .B2 (n_2994));
AOI21_X1 i_978 (.ZN (n_3113), .A (n_2984), .B1 (n_2986), .B2 (n_2987));
AOI22_X1 i_977 (.ZN (n_3112), .A1 (n_1041), .A2 (n_3110), .B1 (n_1048), .B2 (n_1043));
INV_X1 i_975 (.ZN (n_3110), .A (n_1040));
XOR2_X1 i_974 (.Z (n_3109), .A (n_3100), .B (n_3108));
XNOR2_X1 i_973 (.ZN (n_3108), .A (n_4123), .B (n_4117));
XNOR2_X1 i_972 (.ZN (n_3100), .A (n_4154), .B (n_4136));
XNOR2_X1 i_971 (.ZN (n_3094), .A (n_3088), .B (n_3093));
XOR2_X1 i_970 (.Z (n_3093), .A (n_3091), .B (n_3092));
AOI22_X1 i_969 (.ZN (n_3092), .A1 (n_2886), .A2 (n_2892), .B1 (n_2878), .B2 (n_2885));
XNOR2_X1 i_968 (.ZN (n_3091), .A (n_3089), .B (n_3090));
AOI22_X1 i_967 (.ZN (n_3090), .A1 (n_2989), .A2 (n_2995), .B1 (n_2982), .B2 (n_2988));
AOI22_X1 i_966 (.ZN (n_3089), .A1 (n_2906), .A2 (n_2912), .B1 (n_2897), .B2 (n_2905));
AOI22_X1 i_965 (.ZN (n_3088), .A1 (n_720), .A2 (n_711), .B1 (n_3086), .B2 (n_3087));
INV_X1 i_964 (.ZN (n_3087), .A (n_721));
INV_X1 i_963 (.ZN (n_3086), .A (n_757));
OAI21_X1 i_962 (.ZN (n_3085), .A (n_3084), .B1 (n_3065), .B2 (n_3083));
NAND2_X1 i_961 (.ZN (n_3084), .A1 (n_3065), .A2 (n_3083));
XOR2_X1 i_960 (.Z (n_3083), .A (n_3067), .B (n_3082));
OAI21_X1 i_959 (.ZN (n_3082), .A (n_3081), .B1 (n_3080), .B2 (n_3077));
NAND2_X1 i_958 (.ZN (n_3081), .A1 (n_3077), .A2 (n_3080));
OAI22_X1 i_957 (.ZN (n_3080), .A1 (n_951), .A2 (n_3078), .B1 (n_3079), .B2 (n_998));
INV_X1 i_956 (.ZN (n_3079), .A (n_952));
INV_X1 i_955 (.ZN (n_3078), .A (n_943));
XNOR2_X1 i_954 (.ZN (n_3077), .A (n_3070), .B (n_3076));
XNOR2_X1 i_953 (.ZN (n_3076), .A (n_4099), .B (n_4098));
XNOR2_X1 i_952 (.ZN (n_3070), .A (n_3068), .B (n_3069));
OAI21_X1 i_951 (.ZN (n_3069), .A (n_1006), .B1 (n_1005), .B2 (n_999));
AOI22_X1 i_950 (.ZN (n_3068), .A1 (n_1020), .A2 (n_1029), .B1 (n_1021), .B2 (n_1024));
AOI22_X1 i_949 (.ZN (n_3067), .A1 (n_1038), .A2 (n_1019), .B1 (n_3066), .B2 (n_1039));
INV_X1 i_948 (.ZN (n_3066), .A (n_1049));
XOR2_X1 i_947 (.Z (n_3065), .A (n_3063), .B (n_3064));
AOI22_X1 i_946 (.ZN (n_3064), .A1 (n_2997), .A2 (n_589), .B1 (n_709), .B2 (n_2996));
AOI22_X1 i_945 (.ZN (n_3063), .A1 (n_1137), .A2 (n_2914), .B1 (n_2913), .B2 (n_2893));
AOI22_X1 i_944 (.ZN (n_3062), .A1 (n_1220), .A2 (n_2918), .B1 (n_2915), .B2 (n_3061));
INV_X1 i_943 (.ZN (n_3061), .A (n_2917));
XOR2_X1 i_942 (.Z (n_3060), .A (n_3057), .B (n_3059));
AOI22_X1 i_941 (.ZN (n_3059), .A1 (n_3058), .A2 (n_3001), .B1 (n_3000), .B2 (n_883));
INV_X1 i_940 (.ZN (n_3058), .A (n_2922));
XNOR2_X1 i_939 (.ZN (n_3057), .A (n_3055), .B (n_3056));
AOI22_X1 i_938 (.ZN (n_3056), .A1 (n_2974), .A2 (n_2999), .B1 (n_2973), .B2 (n_710));
XOR2_X1 i_937 (.Z (n_3055), .A (n_3005), .B (n_3054));
XOR2_X1 i_936 (.Z (n_3054), .A (n_3037), .B (n_3053));
XNOR2_X1 i_935 (.ZN (n_3053), .A (n_3046), .B (n_3052));
XNOR2_X1 i_934 (.ZN (n_3052), .A (n_4335), .B (n_4334));
XOR2_X1 i_933 (.Z (n_3046), .A (n_3041), .B (n_3045));
XNOR2_X1 i_932 (.ZN (n_3045), .A (n_4367), .B (n_3044));
NAND2_X1 i_931 (.ZN (n_3044), .A1 (inputB[10]), .A2 (inputA[27]));
XNOR2_X1 i_930 (.ZN (n_3041), .A (n_4353), .B (n_4351));
XOR2_X1 i_929 (.Z (n_3037), .A (n_3016), .B (n_3036));
OAI21_X1 i_928 (.ZN (n_3036), .A (n_3035), .B1 (n_3028), .B2 (n_3034));
NAND2_X1 i_927 (.ZN (n_3035), .A1 (n_3028), .A2 (n_3034));
XNOR2_X1 i_926 (.ZN (n_3034), .A (n_4051), .B (n_4050));
XOR2_X1 i_925 (.Z (n_3028), .A (n_3021), .B (n_3027));
XNOR2_X1 i_924 (.ZN (n_3027), .A (n_4319), .B (n_4028));
XNOR2_X1 i_923 (.ZN (n_3021), .A (n_4345), .B (n_4344));
XOR2_X1 i_922 (.Z (n_3016), .A (n_3006), .B (n_3015));
XOR2_X1 i_921 (.Z (n_3015), .A (n_3010), .B (n_3014));
XOR2_X1 i_920 (.Z (n_3014), .A (n_4058), .B (n_4057));
XOR2_X1 i_919 (.Z (n_3010), .A (n_4062), .B (n_2983));
AOI22_X1 i_918 (.ZN (n_3006), .A1 (n_719), .A2 (n_714), .B1 (n_715), .B2 (n_717));
AOI22_X1 i_917 (.ZN (n_3005), .A1 (n_940), .A2 (n_884), .B1 (n_1017), .B2 (n_942));
OAI21_X1 i_916 (.ZN (n_3004), .A (n_2869), .B1 (n_2867), .B2 (n_3003));
XNOR2_X1 i_3040 (.ZN (result[36]), .A (n_2870), .B (n_3003));
XNOR2_X1 i_915 (.ZN (n_3003), .A (n_2921), .B (n_3002));
XNOR2_X1 i_914 (.ZN (n_3002), .A (n_2922), .B (n_3001));
XOR2_X1 i_913 (.Z (n_3001), .A (n_883), .B (n_3000));
XNOR2_X1 i_912 (.ZN (n_3000), .A (n_2974), .B (n_2999));
XNOR2_X1 i_911 (.ZN (n_2999), .A (n_2997), .B (n_589));
XOR2_X1 i_910 (.Z (n_2997), .A (n_709), .B (n_2996));
XOR2_X1 i_909 (.Z (n_2996), .A (n_2989), .B (n_2995));
XOR2_X1 i_908 (.Z (n_2995), .A (n_2993), .B (n_2994));
NOR2_X1 i_907 (.ZN (n_2994), .A1 (n_1551), .A2 (n_127));
NOR2_X1 i_906 (.ZN (n_2993), .A1 (n_2991), .A2 (n_2992));
AOI22_X1 i_905 (.ZN (n_2992), .A1 (inputA[10]), .A2 (inputB[26]), .B1 (inputA[9]), .B2 (inputB[27]));
NOR2_X1 i_904 (.ZN (n_2991), .A1 (n_763), .A2 (n_4060));
XOR2_X1 i_903 (.Z (n_2989), .A (n_2982), .B (n_2988));
XOR2_X1 i_902 (.Z (n_2988), .A (n_2986), .B (n_2987));
NAND2_X1 i_901 (.ZN (n_2987), .A1 (inputA[5]), .A2 (inputB[31]));
NOR2_X1 i_900 (.ZN (n_2986), .A1 (n_2984), .A2 (n_2985));
AOI22_X1 i_899 (.ZN (n_2985), .A1 (inputA[6]), .A2 (inputB[30]), .B1 (inputA[7]), .B2 (inputB[29]));
NOR2_X1 i_898 (.ZN (n_2984), .A1 (n_767), .A2 (n_2983));
NAND2_X1 i_897 (.ZN (n_2983), .A1 (inputA[7]), .A2 (inputB[30]));
XOR2_X1 i_896 (.Z (n_2982), .A (n_4157), .B (n_2981));
NAND2_X1 i_895 (.ZN (n_2981), .A1 (inputA[11]), .A2 (inputB[25]));
XOR2_X1 i_894 (.Z (n_2974), .A (n_710), .B (n_2973));
AOI22_X1 i_893 (.ZN (n_2973), .A1 (n_2972), .A2 (n_1355), .B1 (n_1357), .B2 (n_1359));
INV_X1 i_892 (.ZN (n_2972), .A (n_1361));
AOI22_X1 i_891 (.ZN (n_2922), .A1 (n_1552), .A2 (n_2779), .B1 (n_1350), .B2 (n_2778));
OAI21_X1 i_890 (.ZN (n_2921), .A (n_2920), .B1 (n_2872), .B2 (n_2919));
NAND2_X1 i_889 (.ZN (n_2920), .A1 (n_2872), .A2 (n_2919));
XNOR2_X1 i_888 (.ZN (n_2919), .A (n_1220), .B (n_2918));
XNOR2_X1 i_887 (.ZN (n_2918), .A (n_2915), .B (n_2917));
AOI22_X1 i_886 (.ZN (n_2917), .A1 (n_2853), .A2 (n_2916), .B1 (n_2832), .B2 (n_2852));
INV_X1 i_885 (.ZN (n_2916), .A (n_2854));
XOR2_X1 i_884 (.Z (n_2915), .A (n_1137), .B (n_2914));
XOR2_X1 i_883 (.Z (n_2914), .A (n_2893), .B (n_2913));
XNOR2_X1 i_882 (.ZN (n_2913), .A (n_2906), .B (n_2912));
XNOR2_X1 i_881 (.ZN (n_2912), .A (n_4150), .B (n_4149));
XOR2_X1 i_880 (.Z (n_2906), .A (n_2897), .B (n_2905));
OAI21_X1 i_879 (.ZN (n_2905), .A (n_4159), .B1 (n_4160), .B2 (n_4163));
AOI22_X1 i_878 (.ZN (n_50), .A1 (inputA[17]), .A2 (inputB[19]), .B1 (inputB[18]), .B2 (inputA[18]));
XNOR2_X1 i_877 (.ZN (n_2897), .A (n_4119), .B (n_4118));
XNOR2_X1 i_876 (.ZN (n_2893), .A (n_2886), .B (n_2892));
XNOR2_X1 i_875 (.ZN (n_2892), .A (n_4129), .B (n_4128));
XOR2_X1 i_874 (.Z (n_2886), .A (n_2878), .B (n_2885));
OAI21_X1 i_873 (.ZN (n_2885), .A (n_4135), .B1 (n_48), .B2 (n_49));
INV_X1 i_872 (.ZN (n_49), .A (n_1016));
NOR2_X1 i_871 (.ZN (n_48), .A1 (n_4133), .A2 (n_2881));
AOI22_X1 i_870 (.ZN (n_2881), .A1 (inputB[11]), .A2 (inputA[25]), .B1 (inputB[12]), .B2 (inputA[24]));
XNOR2_X1 i_869 (.ZN (n_2878), .A (n_4109), .B (n_756));
AOI22_X1 i_868 (.ZN (n_2872), .A1 (n_2856), .A2 (n_2871), .B1 (n_2827), .B2 (n_2855));
INV_X1 i_867 (.ZN (n_2871), .A (n_2858));
NAND2_X1 i_2906 (.ZN (n_2870), .A1 (n_2868), .A2 (n_2869));
NAND2_X1 i_866 (.ZN (n_2869), .A1 (n_2864), .A2 (n_2866));
INV_X1 i_2904 (.ZN (n_2868), .A (n_2867));
NOR2_X1 i_865 (.ZN (n_2867), .A1 (n_2864), .A2 (n_2866));
AOI21_X1 i_864 (.ZN (n_2866), .A (n_2865), .B1 (n_2737), .B2 (n_2780));
INV_X1 i_863 (.ZN (n_2865), .A (n_2860));
OAI22_X1 i_862 (.ZN (n_2864), .A1 (n_2735), .A2 (n_2862), .B1 (n_2736), .B2 (n_2863));
INV_X1 i_861 (.ZN (n_2863), .A (n_2861));
XNOR2_X1 i_2898 (.ZN (result[35]), .A (n_2735), .B (n_2862));
XOR2_X1 i_860 (.Z (n_2862), .A (n_2736), .B (n_2861));
OAI21_X1 i_859 (.ZN (n_2861), .A (n_2860), .B1 (n_2781), .B2 (n_2859));
NAND2_X1 i_858 (.ZN (n_2860), .A1 (n_2781), .A2 (n_2859));
XNOR2_X1 i_857 (.ZN (n_2859), .A (n_2856), .B (n_2858));
AOI22_X1 i_856 (.ZN (n_2858), .A1 (n_2722), .A2 (n_2857), .B1 (n_2663), .B2 (n_2721));
INV_X1 i_855 (.ZN (n_2857), .A (n_2724));
XOR2_X1 i_854 (.Z (n_2856), .A (n_2827), .B (n_2855));
XNOR2_X1 i_853 (.ZN (n_2855), .A (n_2853), .B (n_2854));
AOI22_X1 i_852 (.ZN (n_2854), .A1 (n_2682), .A2 (n_2720), .B1 (n_2699), .B2 (n_2719));
XOR2_X1 i_851 (.Z (n_2853), .A (n_2832), .B (n_2852));
XNOR2_X1 i_850 (.ZN (n_2852), .A (n_648), .B (n_590));
XOR2_X1 i_849 (.Z (n_2832), .A (n_703), .B (n_707));
XNOR2_X1 i_848 (.ZN (n_2827), .A (n_1222), .B (n_1221));
XOR2_X1 i_847 (.Z (n_2781), .A (n_2737), .B (n_2780));
XOR2_X1 i_846 (.Z (n_2780), .A (n_1552), .B (n_2779));
XOR2_X1 i_845 (.Z (n_2779), .A (n_1350), .B (n_2778));
AOI22_X1 i_844 (.ZN (n_2778), .A1 (n_2638), .A2 (n_2639), .B1 (n_2637), .B2 (n_2631));
OAI21_X1 i_843 (.ZN (n_2737), .A (n_2641), .B1 (n_2642), .B2 (n_2643));
AOI22_X1 i_842 (.ZN (n_2736), .A1 (n_2726), .A2 (n_2728), .B1 (n_2644), .B2 (n_2725));
AOI21_X1 i_841 (.ZN (n_2735), .A (n_2733), .B1 (n_2596), .B2 (n_2731));
XNOR2_X1 i_840 (.ZN (result[34]), .A (n_2596), .B (n_2734));
NOR2_X1 i_839 (.ZN (n_2734), .A1 (n_2732), .A2 (n_2733));
NOR2_X1 i_838 (.ZN (n_2733), .A1 (n_2729), .A2 (n_2730));
INV_X1 i_837 (.ZN (n_2732), .A (n_2731));
NAND2_X1 i_836 (.ZN (n_2731), .A1 (n_2729), .A2 (n_2730));
OAI22_X1 i_835 (.ZN (n_2730), .A1 (n_2572), .A2 (n_2592), .B1 (n_2571), .B2 (n_2568));
XNOR2_X1 i_834 (.ZN (n_2729), .A (n_2726), .B (n_2728));
AOI22_X1 i_833 (.ZN (n_2728), .A1 (n_3453), .A2 (n_2591), .B1 (n_2727), .B2 (n_3294));
INV_X1 i_832 (.ZN (n_2727), .A (n_2575));
XOR2_X1 i_831 (.Z (n_2726), .A (n_2644), .B (n_2725));
XOR2_X1 i_830 (.Z (n_2725), .A (n_2722), .B (n_2724));
AOI22_X1 i_829 (.ZN (n_2724), .A1 (n_3295), .A2 (n_3400), .B1 (n_2723), .B2 (n_3407));
INV_X1 i_828 (.ZN (n_2723), .A (n_3408));
XOR2_X1 i_827 (.Z (n_2722), .A (n_2663), .B (n_2721));
XOR2_X1 i_826 (.Z (n_2721), .A (n_2682), .B (n_2720));
XOR2_X1 i_825 (.Z (n_2720), .A (n_2699), .B (n_2719));
XNOR2_X1 i_824 (.ZN (n_2719), .A (n_674), .B (n_675));
XNOR2_X1 i_823 (.ZN (n_2699), .A (n_680), .B (n_681));
XNOR2_X1 i_822 (.ZN (n_2682), .A (n_701), .B (n_702));
XOR2_X1 i_821 (.Z (n_2663), .A (n_1312), .B (n_1225));
XNOR2_X1 i_820 (.ZN (n_2644), .A (n_2642), .B (n_2643));
AOI22_X1 i_819 (.ZN (n_2643), .A1 (n_2538), .A2 (n_2567), .B1 (n_2474), .B2 (n_2537));
OAI21_X1 i_818 (.ZN (n_2642), .A (n_2641), .B1 (n_2614), .B2 (n_2640));
NAND2_X1 i_817 (.ZN (n_2641), .A1 (n_2614), .A2 (n_2640));
XNOR2_X1 i_816 (.ZN (n_2640), .A (n_2638), .B (n_2639));
OAI21_X1 i_815 (.ZN (n_2639), .A (n_2515), .B1 (n_2516), .B2 (n_2536));
XOR2_X1 i_814 (.Z (n_2638), .A (n_2631), .B (n_2637));
XOR2_X1 i_813 (.Z (n_2637), .A (n_1139), .B (n_1152));
XOR2_X1 i_812 (.Z (n_2631), .A (n_899), .B (n_892));
XNOR2_X1 i_811 (.ZN (n_2614), .A (n_1649), .B (n_1553));
OAI21_X1 i_810 (.ZN (n_2596), .A (n_2594), .B1 (n_2595), .B2 (n_2449));
INV_X1 i_809 (.ZN (n_2595), .A (n_2446));
OAI21_X1 i_808 (.ZN (result[33]), .A (n_2594), .B1 (n_2450), .B2 (n_2593));
NAND2_X1 i_807 (.ZN (n_2594), .A1 (n_2450), .A2 (n_2593));
XNOR2_X1 i_806 (.ZN (n_2593), .A (n_2572), .B (n_2592));
XNOR2_X1 i_805 (.ZN (n_2592), .A (n_3453), .B (n_2591));
XNOR2_X1 i_804 (.ZN (n_2591), .A (n_2575), .B (n_3294));
AOI22_X1 i_803 (.ZN (n_2575), .A1 (n_2334), .A2 (n_2386), .B1 (n_2333), .B2 (n_2332));
XNOR2_X1 i_802 (.ZN (n_2572), .A (n_2568), .B (n_2571));
AOI22_X1 i_801 (.ZN (n_2571), .A1 (n_2569), .A2 (n_2390), .B1 (n_2387), .B2 (n_2570));
INV_X1 i_800 (.ZN (n_2570), .A (n_2389));
INV_X1 i_799 (.ZN (n_2569), .A (n_2311));
XNOR2_X1 i_798 (.ZN (n_2568), .A (n_2538), .B (n_2567));
XOR2_X1 i_797 (.Z (n_2567), .A (n_1559), .B (n_1554));
XOR2_X1 i_796 (.Z (n_2538), .A (n_2474), .B (n_2537));
XNOR2_X1 i_795 (.ZN (n_2537), .A (n_2516), .B (n_2536));
XNOR2_X1 i_794 (.ZN (n_2536), .A (n_1143), .B (n_1142));
OAI21_X1 i_793 (.ZN (n_2516), .A (n_2515), .B1 (n_2490), .B2 (n_2514));
NAND2_X1 i_792 (.ZN (n_2515), .A1 (n_2490), .A2 (n_2514));
OAI21_X1 i_791 (.ZN (n_2514), .A (n_1146), .B1 (n_1148), .B2 (n_1147));
AOI22_X1 i_2531 (.ZN (n_47), .A1 (inputA[14]), .A2 (inputB[19]), .B1 (inputA[15]), .B2 (inputB[18]));
XOR2_X1 i_790 (.Z (n_2490), .A (n_895), .B (n_893));
XNOR2_X1 i_789 (.ZN (n_2474), .A (n_1711), .B (n_1653));
XNOR2_X1 i_788 (.ZN (n_2450), .A (n_2446), .B (n_2449));
AOI22_X1 i_787 (.ZN (n_2449), .A1 (n_2443), .A2 (n_2444), .B1 (n_2391), .B2 (n_2442));
OAI21_X1 i_786 (.ZN (result[32]), .A (n_2447), .B1 (n_2305), .B2 (n_2448));
INV_X1 i_785 (.ZN (n_2448), .A (n_2445));
OAI21_X1 i_784 (.ZN (n_2447), .A (n_2446), .B1 (n_2309), .B2 (n_2445));
AOI21_X1 i_783 (.ZN (n_2446), .A (n_2306), .B1 (n_2309), .B2 (n_2445));
XNOR2_X1 i_782 (.ZN (n_2445), .A (n_2443), .B (n_2444));
OAI21_X1 i_781 (.ZN (n_2444), .A (n_2297), .B1 (n_2211), .B2 (n_2298));
XOR2_X1 i_780 (.Z (n_2443), .A (n_2391), .B (n_2442));
XOR2_X1 i_779 (.Z (n_2442), .A (n_3455), .B (n_3454));
INV_X1 i_778 (.ZN (n_41), .A (n_1514));
INV_X1 i_777 (.ZN (n_40), .A (n_833));
XOR2_X1 i_776 (.Z (n_2391), .A (n_2311), .B (n_2390));
XNOR2_X1 i_775 (.ZN (n_2390), .A (n_2387), .B (n_2389));
AOI22_X1 i_774 (.ZN (n_2389), .A1 (n_2294), .A2 (n_2388), .B1 (n_2256), .B2 (n_2293));
INV_X1 i_773 (.ZN (n_2388), .A (n_2295));
XOR2_X1 i_772 (.Z (n_2387), .A (n_2334), .B (n_2386));
XOR2_X1 i_771 (.Z (n_2386), .A (n_1719), .B (n_1718));
XOR2_X1 i_770 (.Z (n_2334), .A (n_2332), .B (n_2333));
AOI22_X1 i_769 (.ZN (n_2333), .A1 (n_3235), .A2 (n_3234), .B1 (n_3291), .B2 (n_3236));
XOR2_X1 i_768 (.Z (n_2332), .A (n_1661), .B (n_1660));
AOI22_X1 i_767 (.ZN (n_39), .A1 (inputA[3]), .A2 (inputB[29]), .B1 (inputA[4]), .B2 (inputB[28]));
AOI22_X1 i_766 (.ZN (n_2311), .A1 (n_2209), .A2 (n_2310), .B1 (n_2177), .B2 (n_3233));
INV_X1 i_765 (.ZN (n_2310), .A (n_2210));
NAND3_X1 i_764 (.ZN (n_2309), .A1 (n_2308), .A2 (n_2301), .A3 (n_2304));
OAI21_X1 i_763 (.ZN (n_2308), .A (n_2307), .B1 (n_2160), .B2 (n_2303));
INV_X1 i_762 (.ZN (n_2307), .A (n_2302));
INV_X1 i_761 (.ZN (n_2306), .A (n_2305));
OR2_X1 i_760 (.ZN (n_2305), .A1 (n_2304), .A2 (n_2301));
OR2_X1 i_759 (.ZN (n_2304), .A1 (n_2028), .A2 (n_2158));
XNOR2_X1 i_758 (.ZN (result[31]), .A (n_2160), .B (n_2303));
XNOR2_X1 i_757 (.ZN (n_2303), .A (n_2158), .B (n_2302));
OAI21_X1 i_756 (.ZN (n_2302), .A (n_2301), .B1 (n_2299), .B2 (n_2300));
NAND2_X1 i_755 (.ZN (n_2301), .A1 (n_2299), .A2 (n_2300));
AOI22_X1 i_754 (.ZN (n_2300), .A1 (n_2089), .A2 (n_2156), .B1 (n_2033), .B2 (n_2088));
XNOR2_X1 i_753 (.ZN (n_2299), .A (n_2211), .B (n_2298));
OAI21_X1 i_752 (.ZN (n_2298), .A (n_2297), .B1 (n_2213), .B2 (n_2296));
NAND2_X1 i_751 (.ZN (n_2297), .A1 (n_2213), .A2 (n_2296));
XOR2_X1 i_750 (.Z (n_2296), .A (n_2294), .B (n_2295));
AOI22_X1 i_749 (.ZN (n_2295), .A1 (n_2145), .A2 (n_2150), .B1 (n_2142), .B2 (n_2144));
XOR2_X1 i_748 (.Z (n_2294), .A (n_2256), .B (n_2293));
XNOR2_X1 i_747 (.ZN (n_2293), .A (n_3348), .B (n_3327));
AOI22_X1 i_746 (.ZN (n_38), .A1 (inputA[10]), .A2 (inputB[21]), .B1 (inputA[9]), .B2 (inputB[22]));
OAI22_X1 i_2305 (.ZN (n_37), .A1 (n_529), .A2 (n_400), .B1 (n_530), .B2 (n_881));
XOR2_X1 i_745 (.Z (n_2256), .A (n_3300), .B (n_3297));
AOI22_X1 i_744 (.ZN (n_35), .A1 (inputB[15]), .A2 (inputA[16]), .B1 (inputB[14]), .B2 (inputA[17]));
NOR2_X1 i_743 (.ZN (n_34), .A1 (n_1471), .A2 (n_853));
AOI22_X1 i_742 (.ZN (n_2213), .A1 (n_2152), .A2 (n_2212), .B1 (n_2123), .B2 (n_2151));
INV_X1 i_741 (.ZN (n_2212), .A (n_2155));
XNOR2_X1 i_740 (.ZN (n_2211), .A (n_2209), .B (n_2210));
AOI22_X1 i_739 (.ZN (n_2210), .A1 (n_2087), .A2 (n_2085), .B1 (n_2034), .B2 (n_2084));
XOR2_X1 i_738 (.Z (n_2209), .A (n_2177), .B (n_3233));
XNOR2_X1 i_737 (.ZN (n_2177), .A (n_3467), .B (n_3459));
OAI21_X1 i_736 (.ZN (n_2160), .A (n_2028), .B1 (n_2027), .B2 (n_2159));
XNOR2_X1 i_735 (.ZN (result[30]), .A (n_2030), .B (n_2159));
OAI21_X1 i_734 (.ZN (n_2159), .A (n_2158), .B1 (n_2032), .B2 (n_2157));
NAND2_X1 i_733 (.ZN (n_2158), .A1 (n_2032), .A2 (n_2157));
XNOR2_X1 i_732 (.ZN (n_2157), .A (n_2089), .B (n_2156));
XOR2_X1 i_731 (.Z (n_2156), .A (n_2152), .B (n_2155));
AOI22_X1 i_730 (.ZN (n_2155), .A1 (n_2153), .A2 (n_2019), .B1 (n_2154), .B2 (n_2018));
INV_X1 i_729 (.ZN (n_2154), .A (n_1959));
INV_X1 i_728 (.ZN (n_2153), .A (n_1958));
XOR2_X1 i_727 (.Z (n_2152), .A (n_2123), .B (n_2151));
XOR2_X1 i_726 (.Z (n_2151), .A (n_2145), .B (n_2150));
XNOR2_X1 i_725 (.ZN (n_2150), .A (n_3323), .B (n_3301));
XOR2_X1 i_724 (.Z (n_2145), .A (n_2142), .B (n_2144));
AOI22_X1 i_723 (.ZN (n_2144), .A1 (n_1997), .A2 (n_2143), .B1 (n_1996), .B2 (n_1977));
INV_X1 i_722 (.ZN (n_2143), .A (n_2017));
XNOR2_X1 i_721 (.ZN (n_2142), .A (n_3353), .B (n_3349));
INV_X1 i_2164 (.ZN (n_33), .A (n_3253));
XOR2_X1 i_720 (.Z (n_2123), .A (n_3469), .B (n_3468));
INV_X1 i_2127 (.ZN (n_32), .A (n_3138));
XOR2_X1 i_719 (.Z (n_2089), .A (n_2033), .B (n_2088));
XNOR2_X1 i_718 (.ZN (n_2088), .A (n_2085), .B (n_2087));
AOI22_X1 i_717 (.ZN (n_2087), .A1 (n_1906), .A2 (n_1920), .B1 (n_2086), .B2 (n_3072));
INV_X1 i_716 (.ZN (n_2086), .A (n_3179));
XOR2_X1 i_715 (.Z (n_2085), .A (n_2034), .B (n_2084));
XNOR2_X1 i_714 (.ZN (n_2084), .A (n_3464), .B (n_3463));
AOI22_X1 i_713 (.ZN (n_2034), .A1 (n_1943), .A2 (n_1949), .B1 (n_3008), .B2 (n_1942));
AOI22_X1 i_712 (.ZN (n_2033), .A1 (n_1951), .A2 (n_1953), .B1 (n_1921), .B2 (n_1950));
OAI21_X1 i_711 (.ZN (n_2032), .A (n_2021), .B1 (n_2031), .B2 (n_1954));
INV_X1 i_710 (.ZN (n_2031), .A (n_1955));
NOR2_X1 i_709 (.ZN (n_2030), .A1 (n_2027), .A2 (n_2029));
INV_X1 i_708 (.ZN (n_2029), .A (n_2028));
OR3_X1 i_707 (.ZN (n_2028), .A1 (n_1884), .A2 (n_2024), .A3 (n_2022));
AOI21_X1 i_706 (.ZN (n_2027), .A (n_2025), .B1 (n_1883), .B2 (n_2026));
XNOR2_X1 i_705 (.ZN (result[29]), .A (n_1885), .B (n_2026));
AOI21_X1 i_704 (.ZN (n_2026), .A (n_2025), .B1 (n_2024), .B2 (n_2022));
NOR2_X1 i_703 (.ZN (n_2025), .A1 (n_2022), .A2 (n_2024));
AOI22_X1 i_702 (.ZN (n_2024), .A1 (n_1818), .A2 (n_1875), .B1 (n_2023), .B2 (n_1817));
INV_X1 i_701 (.ZN (n_2023), .A (n_1761));
OAI21_X1 i_700 (.ZN (n_2022), .A (n_2021), .B1 (n_1956), .B2 (n_2020));
NAND2_X1 i_699 (.ZN (n_2021), .A1 (n_1956), .A2 (n_2020));
XNOR2_X1 i_698 (.ZN (n_2020), .A (n_1958), .B (n_2019));
XNOR2_X1 i_697 (.ZN (n_2019), .A (n_1959), .B (n_2018));
XOR2_X1 i_696 (.Z (n_2018), .A (n_1997), .B (n_2017));
OAI21_X1 i_695 (.ZN (n_2017), .A (n_3256), .B1 (n_3268), .B2 (n_3273));
XOR2_X1 i_694 (.Z (n_1997), .A (n_1977), .B (n_1996));
XOR2_X1 i_693 (.Z (n_1996), .A (n_3418), .B (n_3417));
AOI22_X1 i_2015 (.ZN (n_31), .A1 (inputA[7]), .A2 (inputB[22]), .B1 (inputA[6]), .B2 (inputB[23]));
NAND2_X1 i_692 (.ZN (n_30), .A1 (inputA[9]), .A2 (inputB[20]));
NAND2_X1 i_691 (.ZN (n_29), .A1 (n_1979), .A2 (n_28));
NAND4_X1 i_690 (.ZN (n_28), .A1 (inputA[10]), .A2 (inputA[11]), .A3 (inputB[18]), .A4 (inputB[19]));
OAI22_X1 i_689 (.ZN (n_1979), .A1 (n_4162), .A2 (n_314), .B1 (n_1136), .B2 (n_400));
XOR2_X1 i_688 (.Z (n_1977), .A (n_3247), .B (n_3246));
AOI22_X1 i_2003 (.ZN (n_27), .A1 (inputB[13]), .A2 (inputA[16]), .B1 (inputA[15]), .B2 (inputB[14]));
NOR2_X1 i_2002 (.ZN (n_26), .A1 (n_3168), .A2 (n_1471));
AOI22_X1 i_687 (.ZN (n_1959), .A1 (n_1849), .A2 (n_1851), .B1 (n_1830), .B2 (n_1848));
AOI22_X1 i_686 (.ZN (n_1958), .A1 (n_1872), .A2 (n_1957), .B1 (n_1855), .B2 (n_1871));
INV_X1 i_685 (.ZN (n_1957), .A (n_1873));
XNOR2_X1 i_684 (.ZN (n_1956), .A (n_1954), .B (n_1955));
AOI22_X1 i_683 (.ZN (n_1955), .A1 (n_1854), .A2 (n_1874), .B1 (n_1853), .B2 (n_1852));
XNOR2_X1 i_682 (.ZN (n_1954), .A (n_1951), .B (n_1953));
AOI22_X1 i_681 (.ZN (n_1953), .A1 (n_1815), .A2 (n_1952), .B1 (n_1814), .B2 (n_1776));
INV_X1 i_680 (.ZN (n_1952), .A (n_1816));
XOR2_X1 i_679 (.Z (n_1951), .A (n_1921), .B (n_1950));
XNOR2_X1 i_678 (.ZN (n_1950), .A (n_1943), .B (n_1949));
XOR2_X1 i_677 (.Z (n_1949), .A (n_3312), .B (n_3320));
XOR2_X1 i_676 (.Z (n_1943), .A (n_3008), .B (n_1942));
AOI22_X1 i_675 (.ZN (n_1942), .A1 (n_1775), .A2 (n_1941), .B1 (n_2927), .B2 (n_1774));
INV_X1 i_674 (.ZN (n_1941), .A (n_1762));
INV_X1 i_673 (.ZN (n_25), .A (n_1605));
INV_X1 i_672 (.ZN (n_24), .A (n_1515));
INV_X1 i_671 (.ZN (n_23), .A (n_1604));
XNOR2_X1 i_670 (.ZN (n_1921), .A (n_1906), .B (n_1920));
XNOR2_X1 i_669 (.ZN (n_1920), .A (n_3485), .B (n_3473));
XNOR2_X1 i_668 (.ZN (n_1906), .A (n_3179), .B (n_3072));
NAND2_X1 i_667 (.ZN (n_1885), .A1 (n_1883), .A2 (n_1884));
OR3_X1 i_666 (.ZN (n_1884), .A1 (n_1757), .A2 (n_1753), .A3 (n_1879));
NAND2_X1 i_665 (.ZN (n_1883), .A1 (n_1882), .A2 (n_1879));
OAI21_X1 i_664 (.ZN (n_1882), .A (n_1758), .B1 (n_1759), .B2 (n_1881));
XNOR2_X1 i_663 (.ZN (result[28]), .A (n_1759), .B (n_1881));
AOI21_X1 i_662 (.ZN (n_1881), .A (n_1880), .B1 (n_1878), .B2 (n_1876));
INV_X1 i_661 (.ZN (n_1880), .A (n_1879));
OR2_X1 i_660 (.ZN (n_1879), .A1 (n_1876), .A2 (n_1878));
INV_X1 i_659 (.ZN (n_1878), .A (n_1877));
AOI22_X1 i_658 (.ZN (n_1877), .A1 (n_1749), .A2 (n_1674), .B1 (n_1671), .B2 (n_1673));
XNOR2_X1 i_657 (.ZN (n_1876), .A (n_1818), .B (n_1875));
XNOR2_X1 i_656 (.ZN (n_1875), .A (n_1854), .B (n_1874));
XOR2_X1 i_655 (.Z (n_1874), .A (n_1872), .B (n_1873));
AOI22_X1 i_654 (.ZN (n_1873), .A1 (n_1676), .A2 (n_1713), .B1 (n_1696), .B2 (n_1712));
XOR2_X1 i_653 (.Z (n_1872), .A (n_1855), .B (n_1871));
XOR2_X1 i_652 (.Z (n_1871), .A (n_3477), .B (n_3475));
AOI22_X1 i_651 (.ZN (n_1855), .A1 (n_1632), .A2 (n_1654), .B1 (n_1631), .B2 (n_1630));
XOR2_X1 i_650 (.Z (n_1854), .A (n_1852), .B (n_1853));
AOI22_X1 i_649 (.ZN (n_1853), .A1 (n_1667), .A2 (n_1670), .B1 (n_1655), .B2 (n_1666));
XNOR2_X1 i_648 (.ZN (n_1852), .A (n_1849), .B (n_1851));
AOI22_X1 i_647 (.ZN (n_1851), .A1 (n_1665), .A2 (n_1659), .B1 (n_1850), .B2 (n_1658));
INV_X1 i_646 (.ZN (n_1850), .A (n_1656));
XOR2_X1 i_645 (.Z (n_1849), .A (n_1830), .B (n_1848));
XNOR2_X1 i_644 (.ZN (n_1848), .A (n_3316), .B (n_3315));
XNOR2_X1 i_643 (.ZN (n_1830), .A (n_3496), .B (n_3488));
XNOR2_X1 i_642 (.ZN (n_1818), .A (n_1761), .B (n_1817));
XOR2_X1 i_641 (.Z (n_1817), .A (n_1815), .B (n_1816));
AOI22_X1 i_640 (.ZN (n_1816), .A1 (n_1746), .A2 (n_1747), .B1 (n_1734), .B2 (n_1745));
XOR2_X1 i_639 (.Z (n_1815), .A (n_1776), .B (n_1814));
XOR2_X1 i_638 (.Z (n_1814), .A (n_3182), .B (n_3195));
AOI22_X1 i_1831 (.ZN (n_22), .A1 (inputA[7]), .A2 (inputB[21]), .B1 (inputA[8]), .B2 (inputB[20]));
XOR2_X1 i_637 (.Z (n_1776), .A (n_1762), .B (n_1775));
XOR2_X1 i_636 (.Z (n_1775), .A (n_2927), .B (n_1774));
AOI22_X1 i_635 (.ZN (n_1774), .A1 (n_1691), .A2 (n_1695), .B1 (n_1683), .B2 (n_1690));
AOI22_X1 i_634 (.ZN (n_1762), .A1 (n_1743), .A2 (n_1744), .B1 (n_1742), .B2 (n_1741));
AOI22_X1 i_633 (.ZN (n_1761), .A1 (n_1715), .A2 (n_1748), .B1 (n_1760), .B2 (n_1714));
INV_X1 i_632 (.ZN (n_1760), .A (n_1675));
OAI21_X1 i_631 (.ZN (n_1759), .A (n_1758), .B1 (n_1757), .B2 (n_1753));
NAND2_X1 i_630 (.ZN (n_1758), .A1 (n_1757), .A2 (n_1753));
OAI21_X1 i_629 (.ZN (n_1757), .A (n_1625), .B1 (n_1756), .B2 (n_1755));
INV_X1 i_628 (.ZN (n_1756), .A (n_1626));
XNOR2_X1 i_627 (.ZN (result[27]), .A (n_1627), .B (n_1755));
AOI21_X1 i_626 (.ZN (n_1755), .A (n_1754), .B1 (n_1752), .B2 (n_1750));
INV_X1 i_625 (.ZN (n_1754), .A (n_1753));
OR2_X1 i_624 (.ZN (n_1753), .A1 (n_1750), .A2 (n_1752));
INV_X1 i_623 (.ZN (n_1752), .A (n_1751));
AOI22_X1 i_622 (.ZN (n_1751), .A1 (n_1526), .A2 (n_1613), .B1 (n_1524), .B2 (n_1525));
XOR2_X1 i_621 (.Z (n_1750), .A (n_1674), .B (n_1749));
XNOR2_X1 i_620 (.ZN (n_1749), .A (n_1715), .B (n_1748));
XNOR2_X1 i_619 (.ZN (n_1748), .A (n_1746), .B (n_1747));
AOI22_X1 i_618 (.ZN (n_1747), .A1 (n_1590), .A2 (n_1609), .B1 (n_2697), .B2 (n_1589));
XOR2_X1 i_617 (.Z (n_1746), .A (n_1734), .B (n_1745));
XNOR2_X1 i_616 (.ZN (n_1745), .A (n_1743), .B (n_1744));
AOI22_X1 i_615 (.ZN (n_1744), .A1 (n_1602), .A2 (n_1608), .B1 (n_1596), .B2 (n_1601));
XOR2_X1 i_614 (.Z (n_1743), .A (n_1741), .B (n_1742));
AOI22_X1 i_613 (.ZN (n_1742), .A1 (n_1584), .A2 (n_1588), .B1 (n_1578), .B2 (n_1583));
XNOR2_X1 i_612 (.ZN (n_1741), .A (n_2970), .B (n_2961));
XNOR2_X1 i_611 (.ZN (n_1734), .A (n_3200), .B (n_3199));
XNOR2_X1 i_610 (.ZN (n_1715), .A (n_1675), .B (n_1714));
XOR2_X1 i_609 (.Z (n_1714), .A (n_1676), .B (n_1713));
XOR2_X1 i_608 (.Z (n_1713), .A (n_1696), .B (n_1712));
OAI21_X1 i_607 (.ZN (n_1712), .A (n_3489), .B1 (n_3491), .B2 (n_3490));
NAND2_X1 i_606 (.ZN (n_21), .A1 (inputA[9]), .A2 (inputB[18]));
NAND2_X1 i_605 (.ZN (n_20), .A1 (inputA[11]), .A2 (inputB[16]));
AOI22_X1 i_604 (.ZN (n_19), .A1 (inputA[13]), .A2 (inputB[14]), .B1 (inputA[12]), .B2 (inputB[15]));
XNOR2_X1 i_603 (.ZN (n_1696), .A (n_1691), .B (n_1695));
XNOR2_X1 i_602 (.ZN (n_1695), .A (n_3377), .B (n_3376));
XOR2_X1 i_601 (.Z (n_1691), .A (n_1683), .B (n_1690));
OAI21_X1 i_600 (.ZN (n_1690), .A (n_18), .B1 (n_1687), .B2 (n_1688));
NAND2_X1 i_599 (.ZN (n_18), .A1 (n_1687), .A2 (n_1688));
INV_X1 i_598 (.ZN (n_1688), .A (n_2968));
NOR2_X1 i_597 (.ZN (n_1687), .A1 (n_3381), .A2 (n_1686));
AOI22_X1 i_596 (.ZN (n_1686), .A1 (inputB[6]), .A2 (inputA[21]), .B1 (inputB[5]), .B2 (inputA[22]));
XNOR2_X1 i_595 (.ZN (n_1683), .A (n_2934), .B (n_2933));
AOI22_X1 i_594 (.ZN (n_1676), .A1 (n_1518), .A2 (n_1519), .B1 (n_1505), .B2 (n_1517));
AOI22_X1 i_593 (.ZN (n_1675), .A1 (n_1522), .A2 (n_1523), .B1 (n_1520), .B2 (n_1521));
XOR2_X1 i_592 (.Z (n_1674), .A (n_1671), .B (n_1673));
AOI22_X1 i_591 (.ZN (n_1673), .A1 (n_1611), .A2 (n_1672), .B1 (n_1558), .B2 (n_1610));
INV_X1 i_590 (.ZN (n_1672), .A (n_1612));
XNOR2_X1 i_589 (.ZN (n_1671), .A (n_1667), .B (n_1670));
AOI22_X1 i_588 (.ZN (n_1670), .A1 (n_1534), .A2 (n_1668), .B1 (n_1669), .B2 (n_1533));
INV_X1 i_587 (.ZN (n_1669), .A (n_1528));
INV_X1 i_586 (.ZN (n_1668), .A (n_1557));
XOR2_X1 i_585 (.Z (n_1667), .A (n_1655), .B (n_1666));
XNOR2_X1 i_584 (.ZN (n_1666), .A (n_1659), .B (n_1665));
XNOR2_X1 i_583 (.ZN (n_1665), .A (n_3535), .B (n_3480));
XNOR2_X1 i_582 (.ZN (n_1659), .A (n_1656), .B (n_1658));
AOI22_X1 i_581 (.ZN (n_1658), .A1 (n_1510), .A2 (n_1516), .B1 (n_1507), .B2 (n_1657));
INV_X1 i_580 (.ZN (n_1657), .A (n_1509));
OAI22_X1 i_579 (.ZN (n_1656), .A1 (n_2712), .A2 (n_2698), .B1 (n_2706), .B2 (n_2700));
XNOR2_X1 i_578 (.ZN (n_1655), .A (n_1632), .B (n_1654));
XNOR2_X1 i_577 (.ZN (n_1654), .A (n_3500), .B (n_3499));
XOR2_X1 i_576 (.Z (n_1632), .A (n_1630), .B (n_1631));
OAI21_X1 i_575 (.ZN (n_1631), .A (n_1556), .B1 (n_1548), .B2 (n_1541));
AOI22_X1 i_574 (.ZN (n_1630), .A1 (n_1628), .A2 (n_1532), .B1 (n_1629), .B2 (n_1530));
INV_X1 i_573 (.ZN (n_1629), .A (n_1531));
INV_X1 i_572 (.ZN (n_1628), .A (n_1529));
NAND2_X1 i_571 (.ZN (n_1627), .A1 (n_1625), .A2 (n_1626));
OR3_X1 i_570 (.ZN (n_1626), .A1 (n_1624), .A2 (n_1383), .A3 (n_1618));
OAI211_X1 i_569 (.ZN (n_1625), .A (n_1618), .B (n_1623), .C1 (n_1624), .C2 (n_1620));
INV_X1 i_568 (.ZN (n_1624), .A (n_1504));
INV_X1 i_567 (.ZN (n_1623), .A (n_1621));
XOR2_X1 i_566 (.Z (result[26]), .A (n_1504), .B (n_1622));
NOR2_X1 i_565 (.ZN (n_1622), .A1 (n_1620), .A2 (n_1621));
NOR2_X1 i_564 (.ZN (n_1621), .A1 (n_1619), .A2 (n_1383));
AND2_X1 i_563 (.ZN (n_1620), .A1 (n_1383), .A2 (n_1619));
OAI21_X1 i_562 (.ZN (n_1619), .A (n_1618), .B1 (n_1614), .B2 (n_1617));
NAND2_X1 i_561 (.ZN (n_1618), .A1 (n_1614), .A2 (n_1617));
AOI21_X1 i_560 (.ZN (n_1617), .A (n_1615), .B1 (n_1616), .B2 (n_1406));
INV_X1 i_559 (.ZN (n_1616), .A (n_1386));
INV_X1 i_558 (.ZN (n_1615), .A (n_1497));
XNOR2_X1 i_557 (.ZN (n_1614), .A (n_1526), .B (n_1613));
XOR2_X1 i_556 (.Z (n_1613), .A (n_1611), .B (n_1612));
AOI22_X1 i_555 (.ZN (n_1612), .A1 (n_1387), .A2 (n_1405), .B1 (n_1404), .B2 (n_1403));
XOR2_X1 i_554 (.Z (n_1611), .A (n_1558), .B (n_1610));
XOR2_X1 i_553 (.Z (n_1610), .A (n_1590), .B (n_1609));
XNOR2_X1 i_552 (.ZN (n_1609), .A (n_1602), .B (n_1608));
XNOR2_X1 i_551 (.ZN (n_1608), .A (n_2950), .B (n_2949));
XOR2_X1 i_550 (.Z (n_1602), .A (n_1596), .B (n_1601));
XNOR2_X1 i_549 (.ZN (n_1601), .A (n_2955), .B (n_2954));
XOR2_X1 i_548 (.Z (n_1596), .A (n_2964), .B (n_2963));
XOR2_X1 i_547 (.Z (n_1590), .A (n_2697), .B (n_1589));
XNOR2_X1 i_546 (.ZN (n_1589), .A (n_1584), .B (n_1588));
XNOR2_X1 i_545 (.ZN (n_1588), .A (n_3040), .B (n_1587));
NAND2_X1 i_544 (.ZN (n_1587), .A1 (inputA[6]), .A2 (inputB[20]));
XOR2_X1 i_543 (.Z (n_1584), .A (n_1578), .B (n_1583));
XNOR2_X1 i_542 (.ZN (n_1583), .A (n_3048), .B (n_3047));
XOR2_X1 i_541 (.Z (n_1578), .A (n_2941), .B (n_2940));
XOR2_X1 i_540 (.Z (n_1558), .A (n_1534), .B (n_1557));
OAI21_X1 i_539 (.ZN (n_1557), .A (n_1556), .B1 (n_1549), .B2 (n_1555));
NAND2_X1 i_538 (.ZN (n_1556), .A1 (n_1549), .A2 (n_1555));
XNOR2_X1 i_537 (.ZN (n_1555), .A (n_3218), .B (n_3206));
XOR2_X1 i_536 (.Z (n_1549), .A (n_1541), .B (n_1548));
XOR2_X1 i_535 (.Z (n_1548), .A (n_3540), .B (n_3536));
XOR2_X1 i_534 (.Z (n_1541), .A (n_3507), .B (n_17));
AOI21_X1 i_533 (.ZN (n_17), .A (n_1457), .B1 (n_1459), .B2 (n_1539));
INV_X1 i_532 (.ZN (n_1539), .A (n_3071));
XNOR2_X1 i_531 (.ZN (n_1534), .A (n_1528), .B (n_1533));
XOR2_X1 i_530 (.Z (n_1533), .A (n_1529), .B (n_1532));
XNOR2_X1 i_529 (.ZN (n_1532), .A (n_1530), .B (n_1531));
AOI22_X1 i_528 (.ZN (n_1531), .A1 (n_1449), .A2 (n_1454), .B1 (n_1444), .B2 (n_1448));
OAI21_X1 i_527 (.ZN (n_1530), .A (n_1476), .B1 (n_1468), .B2 (n_1461));
AOI22_X1 i_526 (.ZN (n_1529), .A1 (n_1486), .A2 (n_1491), .B1 (n_1484), .B2 (n_1485));
AOI22_X1 i_525 (.ZN (n_1528), .A1 (n_1388), .A2 (n_1402), .B1 (n_1527), .B2 (n_1401));
INV_X1 i_524 (.ZN (n_1527), .A (n_1390));
XOR2_X1 i_523 (.Z (n_1526), .A (n_1524), .B (n_1525));
OAI21_X1 i_522 (.ZN (n_1525), .A (n_1494), .B1 (n_1495), .B2 (n_2789));
XNOR2_X1 i_521 (.ZN (n_1524), .A (n_1522), .B (n_1523));
AOI22_X1 i_520 (.ZN (n_1523), .A1 (n_2806), .A2 (n_2790), .B1 (n_2851), .B2 (n_2807));
XOR2_X1 i_519 (.Z (n_1522), .A (n_1520), .B (n_1521));
AOI22_X1 i_518 (.ZN (n_1521), .A1 (n_1492), .A2 (n_1478), .B1 (n_1455), .B2 (n_1477));
XNOR2_X1 i_517 (.ZN (n_1520), .A (n_1518), .B (n_1519));
AOI22_X1 i_516 (.ZN (n_1519), .A1 (n_2825), .A2 (n_2808), .B1 (n_2831), .B2 (n_2826));
XOR2_X1 i_515 (.Z (n_1518), .A (n_1505), .B (n_1517));
XNOR2_X1 i_514 (.ZN (n_1517), .A (n_1510), .B (n_1516));
XOR2_X1 i_513 (.Z (n_1516), .A (n_2979), .B (n_2978));
XNOR2_X1 i_512 (.ZN (n_1510), .A (n_1507), .B (n_1509));
AOI22_X1 i_511 (.ZN (n_1509), .A1 (n_1481), .A2 (n_1483), .B1 (n_1479), .B2 (n_1508));
INV_X1 i_510 (.ZN (n_1508), .A (n_3007));
OAI22_X1 i_509 (.ZN (n_1507), .A1 (n_2814), .A2 (n_2809), .B1 (n_2819), .B2 (n_1506));
INV_X1 i_508 (.ZN (n_1506), .A (n_2815));
AOI22_X1 i_507 (.ZN (n_1505), .A1 (n_2804), .A2 (n_2791), .B1 (n_2792), .B2 (n_2798));
AOI21_X1 i_506 (.ZN (n_1504), .A (n_1503), .B1 (n_1380), .B2 (n_1501));
INV_X1 i_505 (.ZN (n_1503), .A (n_1500));
XOR2_X1 i_504 (.Z (result[25]), .A (n_1380), .B (n_1502));
NAND2_X1 i_503 (.ZN (n_1502), .A1 (n_1500), .A2 (n_1501));
OR2_X1 i_502 (.ZN (n_1501), .A1 (n_1385), .A2 (n_1499));
NAND2_X1 i_501 (.ZN (n_1500), .A1 (n_1385), .A2 (n_1499));
INV_X1 i_500 (.ZN (n_1499), .A (n_1498));
OAI21_X1 i_499 (.ZN (n_1498), .A (n_1497), .B1 (n_1407), .B2 (n_1496));
NAND2_X1 i_498 (.ZN (n_1497), .A1 (n_1407), .A2 (n_1496));
XOR2_X1 i_497 (.Z (n_1496), .A (n_2789), .B (n_1495));
OAI21_X1 i_496 (.ZN (n_1495), .A (n_1494), .B1 (n_1438), .B2 (n_1493));
NAND2_X1 i_495 (.ZN (n_1494), .A1 (n_1438), .A2 (n_1493));
XOR2_X1 i_494 (.Z (n_1493), .A (n_1478), .B (n_1492));
XNOR2_X1 i_493 (.ZN (n_1492), .A (n_1486), .B (n_1491));
XOR2_X1 i_492 (.Z (n_1491), .A (n_3562), .B (n_1490));
NAND2_X1 i_491 (.ZN (n_1490), .A1 (inputB[4]), .A2 (inputA[21]));
XOR2_X1 i_490 (.Z (n_1486), .A (n_1484), .B (n_1485));
OAI22_X1 i_489 (.ZN (n_1485), .A1 (n_1365), .A2 (n_1366), .B1 (n_1363), .B2 (n_1364));
XOR2_X1 i_488 (.Z (n_1484), .A (n_1481), .B (n_1483));
NOR2_X1 i_487 (.ZN (n_1483), .A1 (n_63), .A2 (n_585));
XNOR2_X1 i_486 (.ZN (n_1481), .A (n_1479), .B (n_3007));
OAI22_X1 i_485 (.ZN (n_1479), .A1 (n_2924), .A2 (n_2923), .B1 (n_2926), .B2 (n_2925));
XOR2_X1 i_484 (.Z (n_1478), .A (n_1455), .B (n_1477));
OAI21_X1 i_483 (.ZN (n_1477), .A (n_1476), .B1 (n_1469), .B2 (n_1475));
NAND2_X1 i_482 (.ZN (n_1476), .A1 (n_1469), .A2 (n_1475));
XOR2_X1 i_481 (.Z (n_1475), .A (n_3215), .B (n_3214));
XOR2_X1 i_480 (.Z (n_1469), .A (n_1461), .B (n_1468));
OAI21_X1 i_479 (.ZN (n_1468), .A (n_3517), .B1 (n_3518), .B2 (n_3534));
XOR2_X1 i_478 (.Z (n_1461), .A (n_1459), .B (n_3071));
NOR2_X1 i_477 (.ZN (n_1459), .A1 (n_1457), .A2 (n_1458));
AOI22_X1 i_476 (.ZN (n_1458), .A1 (inputA[10]), .A2 (inputB[15]), .B1 (inputA[11]), .B2 (inputB[14]));
NOR2_X1 i_475 (.ZN (n_1457), .A1 (n_2850), .A2 (n_3047));
XNOR2_X1 i_474 (.ZN (n_1455), .A (n_1449), .B (n_1454));
XOR2_X1 i_473 (.Z (n_1454), .A (n_3510), .B (n_3509));
XOR2_X1 i_472 (.Z (n_1449), .A (n_1444), .B (n_1448));
XOR2_X1 i_471 (.Z (n_1448), .A (n_3538), .B (n_3537));
XNOR2_X1 i_470 (.ZN (n_1444), .A (n_3543), .B (n_2959));
AOI22_X1 i_469 (.ZN (n_1438), .A1 (n_1372), .A2 (n_1371), .B1 (n_1437), .B2 (n_1370));
INV_X1 i_468 (.ZN (n_1437), .A (n_1354));
XNOR2_X1 i_467 (.ZN (n_1407), .A (n_1386), .B (n_1406));
XNOR2_X1 i_466 (.ZN (n_1406), .A (n_1387), .B (n_1405));
XOR2_X1 i_465 (.Z (n_1405), .A (n_1403), .B (n_1404));
OAI22_X1 i_464 (.ZN (n_1404), .A1 (n_1279), .A2 (n_1319), .B1 (n_1299), .B2 (n_1318));
XNOR2_X1 i_463 (.ZN (n_1403), .A (n_1388), .B (n_1402));
XNOR2_X1 i_462 (.ZN (n_1402), .A (n_1390), .B (n_1401));
XNOR2_X1 i_461 (.ZN (n_1401), .A (n_1397), .B (n_2714));
NAND2_X1 i_460 (.ZN (n_1397), .A1 (n_2755), .A2 (n_2754));
AOI22_X1 i_459 (.ZN (n_1390), .A1 (n_1368), .A2 (n_1389), .B1 (n_1362), .B2 (n_1367));
INV_X1 i_458 (.ZN (n_1389), .A (n_1369));
AOI22_X1 i_457 (.ZN (n_1388), .A1 (n_1329), .A2 (n_1335), .B1 (n_1323), .B2 (n_1328));
AOI22_X1 i_456 (.ZN (n_1387), .A1 (n_1338), .A2 (n_1351), .B1 (n_1337), .B2 (n_1336));
AOI22_X1 i_455 (.ZN (n_1386), .A1 (n_1321), .A2 (n_1352), .B1 (n_1278), .B2 (n_1320));
AOI22_X1 i_454 (.ZN (n_1385), .A1 (n_1383), .A2 (n_1384), .B1 (n_1353), .B2 (n_1375));
OAI21_X1 i_453 (.ZN (n_1384), .A (n_1381), .B1 (n_1382), .B2 (n_1373));
OR3_X1 i_452 (.ZN (n_1383), .A1 (n_1381), .A2 (n_1382), .A3 (n_1373));
INV_X1 i_451 (.ZN (n_1382), .A (n_1374));
NAND2_X1 i_450 (.ZN (n_1381), .A1 (n_1376), .A2 (n_1377));
AOI21_X1 i_449 (.ZN (n_1380), .A (n_1379), .B1 (n_1274), .B2 (n_1378));
INV_X1 i_448 (.ZN (n_1379), .A (n_1275));
XNOR2_X1 i_447 (.ZN (result[24]), .A (n_1276), .B (n_1378));
XOR2_X1 i_446 (.Z (n_1378), .A (n_1376), .B (n_1377));
OAI21_X1 i_445 (.ZN (n_1377), .A (n_1195), .B1 (n_1196), .B2 (n_1265));
XOR2_X1 i_444 (.Z (n_1376), .A (n_1353), .B (n_1375));
XNOR2_X1 i_443 (.ZN (n_1375), .A (n_1373), .B (n_1374));
OAI21_X1 i_442 (.ZN (n_1374), .A (n_1260), .B1 (n_1261), .B2 (n_1264));
XNOR2_X1 i_441 (.ZN (n_1373), .A (n_1371), .B (n_1372));
AOI22_X1 i_440 (.ZN (n_1372), .A1 (n_1197), .A2 (n_1234), .B1 (n_1233), .B2 (n_1218));
XNOR2_X1 i_439 (.ZN (n_1371), .A (n_1354), .B (n_1370));
XOR2_X1 i_438 (.Z (n_1370), .A (n_1368), .B (n_1369));
AOI22_X1 i_437 (.ZN (n_1369), .A1 (n_1249), .A2 (n_1255), .B1 (n_1248), .B2 (n_1242));
XOR2_X1 i_436 (.Z (n_1368), .A (n_1362), .B (n_1367));
XNOR2_X1 i_435 (.ZN (n_1367), .A (n_1365), .B (n_1366));
NAND2_X1 i_434 (.ZN (n_1366), .A1 (inputB[0]), .A2 (inputA[24]));
XNOR2_X1 i_433 (.ZN (n_1365), .A (n_1363), .B (n_1364));
AOI21_X1 i_432 (.ZN (n_1364), .A (n_2890), .B1 (n_2888), .B2 (n_2887));
AOI21_X1 i_431 (.ZN (n_1363), .A (n_2902), .B1 (n_2900), .B2 (n_2899));
XNOR2_X1 i_430 (.ZN (n_1362), .A (n_2771), .B (n_2765));
AOI22_X1 i_429 (.ZN (n_1354), .A1 (n_1258), .A2 (n_1237), .B1 (n_1257), .B2 (n_1256));
XNOR2_X1 i_428 (.ZN (n_1353), .A (n_1321), .B (n_1352));
XOR2_X1 i_427 (.Z (n_1352), .A (n_1338), .B (n_1351));
XNOR2_X1 i_426 (.ZN (n_1351), .A (n_2903), .B (n_2873));
XOR2_X1 i_425 (.Z (n_1338), .A (n_1336), .B (n_1337));
OAI21_X1 i_424 (.ZN (n_1337), .A (n_2676), .B1 (n_2675), .B2 (n_1176));
XNOR2_X1 i_423 (.ZN (n_1336), .A (n_1329), .B (n_1335));
XNOR2_X1 i_422 (.ZN (n_1335), .A (n_2741), .B (n_2715));
XOR2_X1 i_421 (.Z (n_1329), .A (n_1323), .B (n_1328));
XNOR2_X1 i_420 (.ZN (n_1328), .A (n_2760), .B (n_2759));
AOI22_X1 i_419 (.ZN (n_1323), .A1 (n_1173), .A2 (n_1175), .B1 (n_1322), .B2 (n_1172));
INV_X1 i_418 (.ZN (n_1322), .A (n_1170));
XOR2_X1 i_417 (.Z (n_1321), .A (n_1278), .B (n_1320));
XNOR2_X1 i_416 (.ZN (n_1320), .A (n_1279), .B (n_1319));
XNOR2_X1 i_415 (.ZN (n_1319), .A (n_1299), .B (n_1318));
XOR2_X1 i_414 (.Z (n_1318), .A (n_2794), .B (n_2793));
XOR2_X1 i_413 (.Z (n_1299), .A (n_2800), .B (n_2799));
AOI22_X1 i_412 (.ZN (n_1279), .A1 (n_2635), .A2 (n_1178), .B1 (n_2636), .B2 (n_2657));
AOI22_X1 i_411 (.ZN (n_1278), .A1 (n_1192), .A2 (n_1277), .B1 (n_1177), .B2 (n_1191));
INV_X1 i_410 (.ZN (n_1277), .A (n_1193));
NAND2_X1 i_409 (.ZN (n_1276), .A1 (n_1274), .A2 (n_1275));
OR3_X1 i_408 (.ZN (n_1275), .A1 (n_1271), .A2 (n_1161), .A3 (n_1273));
OAI21_X1 i_407 (.ZN (n_1274), .A (n_1273), .B1 (n_1269), .B2 (n_1267));
NAND2_X1 i_406 (.ZN (n_1273), .A1 (n_1266), .A2 (n_1163));
XOR2_X1 i_405 (.Z (result[23]), .A (n_1267), .B (n_1272));
OAI21_X1 i_404 (.ZN (n_1272), .A (n_1270), .B1 (n_1271), .B2 (n_1161));
INV_X1 i_403 (.ZN (n_1271), .A (n_1071));
INV_X1 i_402 (.ZN (n_1270), .A (n_1269));
NOR2_X1 i_401 (.ZN (n_1269), .A1 (n_1268), .A2 (n_1071));
OAI21_X1 i_400 (.ZN (n_1268), .A (n_1161), .B1 (n_1070), .B2 (n_1162));
XNOR2_X1 i_399 (.ZN (n_1267), .A (n_1163), .B (n_1266));
XOR2_X1 i_398 (.Z (n_1266), .A (n_1196), .B (n_1265));
XNOR2_X1 i_397 (.ZN (n_1265), .A (n_1261), .B (n_1264));
AOI22_X1 i_396 (.ZN (n_1264), .A1 (n_1087), .A2 (n_1262), .B1 (n_1263), .B2 (n_2583));
INV_X1 i_395 (.ZN (n_1263), .A (n_1074));
INV_X1 i_394 (.ZN (n_1262), .A (n_1089));
OAI21_X1 i_393 (.ZN (n_1261), .A (n_1260), .B1 (n_1235), .B2 (n_1259));
NAND2_X1 i_392 (.ZN (n_1260), .A1 (n_1235), .A2 (n_1259));
XOR2_X1 i_391 (.Z (n_1259), .A (n_1237), .B (n_1258));
XOR2_X1 i_390 (.Z (n_1258), .A (n_1256), .B (n_1257));
AOI22_X1 i_389 (.ZN (n_1257), .A1 (n_1115), .A2 (n_1120), .B1 (n_1108), .B2 (n_1114));
XNOR2_X1 i_388 (.ZN (n_1256), .A (n_1249), .B (n_1255));
XOR2_X1 i_387 (.Z (n_1255), .A (n_2717), .B (n_2764));
XOR2_X1 i_386 (.Z (n_1249), .A (n_1242), .B (n_1248));
XNOR2_X1 i_385 (.ZN (n_1248), .A (n_2746), .B (n_2745));
XNOR2_X1 i_384 (.ZN (n_1242), .A (n_2751), .B (n_2750));
AOI22_X1 i_383 (.ZN (n_1237), .A1 (n_2584), .A2 (n_2602), .B1 (n_1236), .B2 (n_2603));
INV_X1 i_382 (.ZN (n_1236), .A (n_2613));
XNOR2_X1 i_381 (.ZN (n_1235), .A (n_1197), .B (n_1234));
XOR2_X1 i_380 (.Z (n_1234), .A (n_1218), .B (n_1233));
XNOR2_X1 i_379 (.ZN (n_1233), .A (n_2894), .B (n_2884));
XOR2_X1 i_378 (.Z (n_1218), .A (n_2880), .B (n_2879));
AOI22_X1 i_377 (.ZN (n_1197), .A1 (n_1105), .A2 (n_1106), .B1 (n_1104), .B2 (n_1092));
OAI21_X1 i_376 (.ZN (n_1196), .A (n_1195), .B1 (n_1164), .B2 (n_1194));
NAND2_X1 i_375 (.ZN (n_1195), .A1 (n_1164), .A2 (n_1194));
XNOR2_X1 i_374 (.ZN (n_1194), .A (n_1192), .B (n_1193));
AOI22_X1 i_373 (.ZN (n_1193), .A1 (n_1121), .A2 (n_1154), .B1 (n_1135), .B2 (n_1153));
XOR2_X1 i_372 (.Z (n_1192), .A (n_1177), .B (n_1191));
XOR2_X1 i_371 (.Z (n_1191), .A (n_1178), .B (n_2635));
AOI22_X1 i_370 (.ZN (n_1178), .A1 (n_1130), .A2 (n_1134), .B1 (n_1125), .B2 (n_1129));
XNOR2_X1 i_369 (.ZN (n_1177), .A (n_2675), .B (n_1176));
XNOR2_X1 i_368 (.ZN (n_1176), .A (n_1173), .B (n_1175));
AOI22_X1 i_367 (.ZN (n_1175), .A1 (n_2606), .A2 (n_2604), .B1 (n_2612), .B2 (n_1174));
INV_X1 i_366 (.ZN (n_1174), .A (n_2607));
XNOR2_X1 i_365 (.ZN (n_1173), .A (n_1170), .B (n_1172));
AOI22_X1 i_364 (.ZN (n_1172), .A1 (n_1111), .A2 (n_1113), .B1 (n_1171), .B2 (n_1110));
INV_X1 i_363 (.ZN (n_1171), .A (n_2740));
OAI22_X1 i_362 (.ZN (n_1170), .A1 (n_1118), .A2 (n_1119), .B1 (n_1116), .B2 (n_1117));
AOI22_X1 i_361 (.ZN (n_1164), .A1 (n_1156), .A2 (n_2582), .B1 (n_1107), .B2 (n_1155));
AOI22_X1 i_360 (.ZN (n_1163), .A1 (n_1091), .A2 (n_1158), .B1 (n_1073), .B2 (n_1090));
XNOR2_X1 i_359 (.ZN (result[22]), .A (n_1072), .B (n_1162));
OAI21_X1 i_358 (.ZN (n_1162), .A (n_1161), .B1 (n_1159), .B2 (n_1160));
NAND2_X1 i_357 (.ZN (n_1161), .A1 (n_1159), .A2 (n_1160));
OAI22_X1 i_356 (.ZN (n_1160), .A1 (n_1063), .A2 (n_1032), .B1 (n_1034), .B2 (n_1062));
XNOR2_X1 i_355 (.ZN (n_1159), .A (n_1091), .B (n_1158));
XOR2_X1 i_354 (.Z (n_1158), .A (n_1156), .B (n_2582));
XOR2_X1 i_353 (.Z (n_1156), .A (n_1107), .B (n_1155));
XNOR2_X1 i_352 (.ZN (n_1155), .A (n_1121), .B (n_1154));
XOR2_X1 i_351 (.Z (n_1154), .A (n_1135), .B (n_1153));
OAI21_X1 i_350 (.ZN (n_1153), .A (n_2679), .B1 (n_2681), .B2 (n_2680));
XNOR2_X1 i_349 (.ZN (n_1135), .A (n_1130), .B (n_1134));
XNOR2_X1 i_348 (.ZN (n_1134), .A (n_2654), .B (n_1133));
NAND2_X1 i_347 (.ZN (n_1133), .A1 (inputA[3]), .A2 (inputB[19]));
XOR2_X1 i_346 (.Z (n_1130), .A (n_1125), .B (n_1129));
XNOR2_X1 i_345 (.ZN (n_1129), .A (n_2647), .B (n_1128));
NAND2_X1 i_344 (.ZN (n_1128), .A1 (inputA[9]), .A2 (inputB[13]));
XNOR2_X1 i_343 (.ZN (n_1125), .A (n_2651), .B (n_2650));
XNOR2_X1 i_342 (.ZN (n_1121), .A (n_1115), .B (n_1120));
XNOR2_X1 i_341 (.ZN (n_1120), .A (n_1118), .B (n_1119));
AOI21_X1 i_340 (.ZN (n_1119), .A (n_984), .B1 (n_986), .B2 (n_987));
XNOR2_X1 i_339 (.ZN (n_1118), .A (n_1116), .B (n_1117));
AOI21_X1 i_338 (.ZN (n_1117), .A (n_2633), .B1 (n_2630), .B2 (n_2629));
AOI21_X1 i_337 (.ZN (n_1116), .A (n_990), .B1 (n_992), .B2 (n_2559));
XOR2_X1 i_336 (.Z (n_1115), .A (n_1108), .B (n_1114));
XNOR2_X1 i_335 (.ZN (n_1114), .A (n_1111), .B (n_1113));
NOR2_X1 i_334 (.ZN (n_1113), .A1 (n_66), .A2 (n_217));
XNOR2_X1 i_333 (.ZN (n_1111), .A (n_1110), .B (n_2740));
NOR2_X1 i_332 (.ZN (n_1110), .A1 (n_67), .A2 (n_414));
AOI22_X1 i_331 (.ZN (n_1108), .A1 (n_978), .A2 (n_981), .B1 (n_979), .B2 (n_980));
XNOR2_X1 i_330 (.ZN (n_1107), .A (n_1105), .B (n_1106));
OAI21_X1 i_329 (.ZN (n_1106), .A (n_995), .B1 (n_988), .B2 (n_993));
XOR2_X1 i_328 (.Z (n_1105), .A (n_1092), .B (n_1104));
XOR2_X1 i_327 (.Z (n_1104), .A (n_2692), .B (n_2685));
AOI22_X1 i_326 (.ZN (n_1092), .A1 (n_2550), .A2 (n_2565), .B1 (n_2543), .B2 (n_2549));
XOR2_X1 i_325 (.Z (n_1091), .A (n_1073), .B (n_1090));
XOR2_X1 i_324 (.Z (n_1090), .A (n_1087), .B (n_1089));
AOI22_X1 i_323 (.ZN (n_1089), .A1 (n_1014), .A2 (n_1030), .B1 (n_1088), .B2 (n_1013));
INV_X1 i_322 (.ZN (n_1088), .A (n_996));
XNOR2_X1 i_321 (.ZN (n_1087), .A (n_1074), .B (n_2583));
AOI22_X1 i_320 (.ZN (n_1074), .A1 (n_2566), .A2 (n_2577), .B1 (n_2574), .B2 (n_2576));
AOI22_X1 i_319 (.ZN (n_1073), .A1 (n_976), .A2 (n_1031), .B1 (n_974), .B2 (n_975));
NOR2_X1 i_318 (.ZN (n_1072), .A1 (n_1070), .A2 (n_1071));
AND2_X1 i_317 (.ZN (n_1071), .A1 (n_1069), .A2 (n_1067));
AOI211_X1 i_316 (.ZN (n_1070), .A (n_1067), .B (n_1069), .C1 (n_971), .C2 (n_1068));
INV_X1 i_315 (.ZN (n_1069), .A (n_972));
XNOR2_X1 i_314 (.ZN (result[21]), .A (n_973), .B (n_1068));
AOI21_X1 i_313 (.ZN (n_1068), .A (n_1067), .B1 (n_1066), .B2 (n_1064));
NOR2_X1 i_312 (.ZN (n_1067), .A1 (n_1064), .A2 (n_1066));
INV_X1 i_311 (.ZN (n_1066), .A (n_1065));
OAI21_X1 i_310 (.ZN (n_1065), .A (n_927), .B1 (n_928), .B2 (n_959));
XNOR2_X1 i_309 (.ZN (n_1064), .A (n_1032), .B (n_1063));
XNOR2_X1 i_308 (.ZN (n_1063), .A (n_1034), .B (n_1062));
XNOR2_X1 i_307 (.ZN (n_1062), .A (n_2578), .B (n_2581));
AOI22_X1 i_306 (.ZN (n_1034), .A1 (n_932), .A2 (n_958), .B1 (n_1033), .B2 (n_931));
INV_X1 i_305 (.ZN (n_1033), .A (n_1795));
XNOR2_X1 i_304 (.ZN (n_1032), .A (n_976), .B (n_1031));
XOR2_X1 i_303 (.Z (n_1031), .A (n_1014), .B (n_1030));
XOR2_X1 i_302 (.Z (n_1030), .A (n_2587), .B (n_2585));
XNOR2_X1 i_301 (.ZN (n_1014), .A (n_996), .B (n_1013));
XNOR2_X1 i_300 (.ZN (n_1013), .A (n_2622), .B (n_2615));
OAI21_X1 i_299 (.ZN (n_996), .A (n_995), .B1 (n_982), .B2 (n_994));
NAND2_X1 i_298 (.ZN (n_995), .A1 (n_982), .A2 (n_994));
XOR2_X1 i_297 (.Z (n_994), .A (n_988), .B (n_993));
XNOR2_X1 i_296 (.ZN (n_993), .A (n_992), .B (n_2559));
NOR2_X1 i_295 (.ZN (n_992), .A1 (n_990), .A2 (n_991));
AOI22_X1 i_294 (.ZN (n_991), .A1 (inputA[1]), .A2 (inputB[20]), .B1 (inputA[0]), .B2 (inputB[21]));
NOR2_X1 i_293 (.ZN (n_990), .A1 (n_2563), .A2 (n_2740));
XNOR2_X1 i_292 (.ZN (n_988), .A (n_986), .B (n_987));
NOR2_X1 i_291 (.ZN (n_987), .A1 (n_1724), .A2 (n_400));
NOR2_X1 i_290 (.ZN (n_986), .A1 (n_984), .A2 (n_985));
AOI22_X1 i_289 (.ZN (n_985), .A1 (inputA[4]), .A2 (inputB[17]), .B1 (inputA[5]), .B2 (inputB[16]));
NOR2_X1 i_288 (.ZN (n_984), .A1 (n_2551), .A2 (n_2656));
XOR2_X1 i_287 (.Z (n_982), .A (n_978), .B (n_981));
XOR2_X1 i_286 (.Z (n_981), .A (n_979), .B (n_980));
OAI21_X1 i_285 (.ZN (n_980), .A (n_2560), .B1 (n_2562), .B2 (n_2563));
OAI22_X1 i_284 (.ZN (n_979), .A1 (n_2555), .A2 (n_2552), .B1 (n_1723), .B2 (n_2551));
OAI22_X1 i_283 (.ZN (n_978), .A1 (n_1902), .A2 (n_1903), .B1 (n_977), .B2 (n_1896));
INV_X1 i_282 (.ZN (n_977), .A (n_1901));
XOR2_X1 i_281 (.Z (n_976), .A (n_974), .B (n_975));
AOI22_X1 i_280 (.ZN (n_975), .A1 (n_956), .A2 (n_1794), .B1 (n_934), .B2 (n_955));
AOI22_X1 i_279 (.ZN (n_974), .A1 (n_1931), .A2 (n_1930), .B1 (n_1965), .B2 (n_1932));
NAND2_X1 i_278 (.ZN (n_973), .A1 (n_971), .A2 (n_972));
NAND2_X1 i_277 (.ZN (n_972), .A1 (n_961), .A2 (n_966));
OAI211_X1 i_276 (.ZN (n_971), .A (n_968), .B (n_962), .C1 (n_969), .C2 (n_970));
INV_X1 i_275 (.ZN (n_970), .A (n_967));
INV_X1 i_274 (.ZN (n_969), .A (n_963));
INV_X1 i_273 (.ZN (n_968), .A (n_966));
XNOR2_X1 i_272 (.ZN (result[20]), .A (n_964), .B (n_967));
AOI21_X1 i_271 (.ZN (n_967), .A (n_966), .B1 (n_870), .B2 (n_965));
NOR2_X1 i_270 (.ZN (n_966), .A1 (n_870), .A2 (n_965));
OAI21_X1 i_269 (.ZN (n_965), .A (n_866), .B1 (n_818), .B2 (n_862));
NAND2_X1 i_268 (.ZN (n_964), .A1 (n_962), .A2 (n_963));
NAND2_X1 i_267 (.ZN (n_963), .A1 (n_875), .A2 (n_960));
INV_X1 i_266 (.ZN (n_962), .A (n_961));
NOR2_X1 i_265 (.ZN (n_961), .A1 (n_875), .A2 (n_960));
XNOR2_X1 i_264 (.ZN (n_960), .A (n_928), .B (n_959));
XNOR2_X1 i_263 (.ZN (n_959), .A (n_932), .B (n_958));
XNOR2_X1 i_262 (.ZN (n_958), .A (n_956), .B (n_1794));
XOR2_X1 i_261 (.Z (n_956), .A (n_934), .B (n_955));
XOR2_X1 i_260 (.Z (n_955), .A (n_947), .B (n_2564));
NAND2_X1 i_259 (.ZN (n_947), .A1 (n_945), .A2 (n_2557));
INV_X1 i_258 (.ZN (n_945), .A (n_2558));
AOI22_X1 i_257 (.ZN (n_934), .A1 (n_789), .A2 (n_933), .B1 (n_783), .B2 (n_788));
INV_X1 i_256 (.ZN (n_933), .A (n_782));
XNOR2_X1 i_255 (.ZN (n_932), .A (n_1795), .B (n_931));
AOI22_X1 i_254 (.ZN (n_931), .A1 (n_861), .A2 (n_820), .B1 (n_840), .B2 (n_930));
INV_X1 i_253 (.ZN (n_930), .A (n_860));
OAI21_X1 i_252 (.ZN (n_928), .A (n_927), .B1 (n_877), .B2 (n_926));
NAND2_X1 i_251 (.ZN (n_927), .A1 (n_877), .A2 (n_926));
XNOR2_X1 i_250 (.ZN (n_926), .A (n_1931), .B (n_1930));
AOI22_X1 i_249 (.ZN (n_877), .A1 (n_791), .A2 (n_817), .B1 (n_876), .B2 (n_790));
INV_X1 i_248 (.ZN (n_876), .A (n_781));
OAI22_X1 i_247 (.ZN (n_875), .A1 (n_780), .A2 (n_872), .B1 (n_873), .B2 (n_874));
INV_X1 i_246 (.ZN (n_874), .A (n_774));
INV_X1 i_245 (.ZN (n_873), .A (n_871));
XNOR2_X1 i_244 (.ZN (result[19]), .A (n_780), .B (n_872));
XNOR2_X1 i_243 (.ZN (n_872), .A (n_871), .B (n_774));
OAI21_X1 i_242 (.ZN (n_871), .A (n_870), .B1 (n_867), .B2 (n_869));
NAND2_X1 i_241 (.ZN (n_870), .A1 (n_867), .A2 (n_869));
AOI22_X1 i_240 (.ZN (n_869), .A1 (n_737), .A2 (n_771), .B1 (n_868), .B2 (n_736));
INV_X1 i_239 (.ZN (n_868), .A (n_696));
OAI21_X1 i_238 (.ZN (n_867), .A (n_866), .B1 (n_863), .B2 (n_2037));
NAND2_X1 i_237 (.ZN (n_866), .A1 (n_863), .A2 (n_2037));
XOR2_X1 i_236 (.Z (n_863), .A (n_818), .B (n_862));
XNOR2_X1 i_235 (.ZN (n_862), .A (n_820), .B (n_861));
XNOR2_X1 i_234 (.ZN (n_861), .A (n_840), .B (n_860));
OAI21_X1 i_233 (.ZN (n_860), .A (n_1998), .B1 (n_2000), .B2 (n_1999));
XNOR2_X1 i_232 (.ZN (n_840), .A (n_2006), .B (n_2004));
AOI22_X1 i_231 (.ZN (n_820), .A1 (n_2039), .A2 (n_2056), .B1 (n_2058), .B2 (n_819));
INV_X1 i_230 (.ZN (n_819), .A (n_2057));
XNOR2_X1 i_229 (.ZN (n_818), .A (n_791), .B (n_817));
XOR2_X1 i_228 (.Z (n_817), .A (n_1797), .B (n_1796));
XNOR2_X1 i_227 (.ZN (n_791), .A (n_781), .B (n_790));
XOR2_X1 i_226 (.Z (n_790), .A (n_782), .B (n_789));
XOR2_X1 i_225 (.Z (n_789), .A (n_783), .B (n_788));
XNOR2_X1 i_224 (.ZN (n_788), .A (n_1983), .B (n_1976));
AOI22_X1 i_223 (.ZN (n_783), .A1 (n_725), .A2 (n_732), .B1 (n_724), .B2 (n_718));
AOI22_X1 i_222 (.ZN (n_782), .A1 (n_2059), .A2 (n_2077), .B1 (n_2082), .B2 (n_2078));
AOI22_X1 i_221 (.ZN (n_781), .A1 (n_735), .A2 (n_734), .B1 (n_713), .B2 (n_733));
AOI21_X1 i_220 (.ZN (n_780), .A (n_778), .B1 (n_694), .B2 (n_779));
INV_X1 i_219 (.ZN (n_779), .A (n_777));
INV_X1 i_218 (.ZN (n_778), .A (n_776));
XOR2_X1 i_217 (.Z (result[18]), .A (n_694), .B (n_777));
OAI21_X1 i_216 (.ZN (n_777), .A (n_776), .B1 (n_625), .B2 (n_775));
NAND2_X1 i_215 (.ZN (n_776), .A1 (n_775), .A2 (n_625));
OAI21_X1 i_214 (.ZN (n_775), .A (n_774), .B1 (n_2410), .B2 (n_772));
NAND2_X1 i_213 (.ZN (n_774), .A1 (n_772), .A2 (n_2410));
XNOR2_X1 i_212 (.ZN (n_772), .A (n_737), .B (n_771));
XNOR2_X1 i_211 (.ZN (n_771), .A (n_2083), .B (n_2038));
XNOR2_X1 i_210 (.ZN (n_737), .A (n_696), .B (n_736));
XOR2_X1 i_209 (.Z (n_736), .A (n_734), .B (n_735));
AOI22_X1 i_208 (.ZN (n_735), .A1 (n_2475), .A2 (n_2459), .B1 (n_2477), .B2 (n_2476));
XOR2_X1 i_207 (.Z (n_734), .A (n_713), .B (n_733));
XOR2_X1 i_206 (.Z (n_733), .A (n_725), .B (n_732));
XNOR2_X1 i_205 (.ZN (n_732), .A (n_1980), .B (n_1978));
XOR2_X1 i_204 (.Z (n_725), .A (n_718), .B (n_724));
XNOR2_X1 i_203 (.ZN (n_724), .A (n_1988), .B (n_1987));
XNOR2_X1 i_202 (.ZN (n_718), .A (n_1992), .B (n_1991));
XOR2_X1 i_201 (.Z (n_713), .A (n_1806), .B (n_1801));
AOI22_X1 i_200 (.ZN (n_696), .A1 (n_2456), .A2 (n_695), .B1 (n_2458), .B2 (n_2457));
INV_X1 i_199 (.ZN (n_695), .A (n_2412));
OAI22_X1 i_198 (.ZN (n_694), .A1 (n_623), .A2 (n_692), .B1 (n_693), .B2 (n_691));
INV_X1 i_197 (.ZN (n_693), .A (n_626));
XNOR2_X1 i_196 (.ZN (result[17]), .A (n_623), .B (n_692));
XOR2_X1 i_195 (.Z (n_692), .A (n_626), .B (n_691));
XOR2_X1 i_194 (.Z (n_691), .A (n_2411), .B (n_2478));
OAI21_X1 i_193 (.ZN (n_626), .A (n_625), .B1 (n_619), .B2 (n_624));
NAND2_X1 i_192 (.ZN (n_625), .A1 (n_624), .A2 (n_619));
AOI22_X1 i_191 (.ZN (n_624), .A1 (n_612), .A2 (n_613), .B1 (n_580), .B2 (n_611));
OAI21_X1 i_190 (.ZN (n_623), .A (n_615), .B1 (n_621), .B2 (n_622));
INV_X1 i_189 (.ZN (n_622), .A (n_620));
INV_X1 i_188 (.ZN (n_621), .A (n_616));
XNOR2_X1 i_187 (.ZN (result[16]), .A (n_617), .B (n_620));
AOI21_X1 i_186 (.ZN (n_620), .A (n_619), .B1 (n_539), .B2 (n_618));
NOR2_X1 i_185 (.ZN (n_619), .A1 (n_539), .A2 (n_618));
AOI22_X1 i_184 (.ZN (n_618), .A1 (n_504), .A2 (n_536), .B1 (n_503), .B2 (n_501));
NAND2_X1 i_183 (.ZN (n_617), .A1 (n_615), .A2 (n_616));
OR2_X1 i_182 (.ZN (n_616), .A1 (n_542), .A2 (n_614));
NAND2_X1 i_181 (.ZN (n_615), .A1 (n_542), .A2 (n_614));
XNOR2_X1 i_180 (.ZN (n_614), .A (n_612), .B (n_613));
AOI22_X1 i_179 (.ZN (n_613), .A1 (n_520), .A2 (n_535), .B1 (n_505), .B2 (n_519));
XOR2_X1 i_178 (.Z (n_612), .A (n_580), .B (n_611));
XOR2_X1 i_177 (.Z (n_611), .A (n_2413), .B (n_2453));
XOR2_X1 i_176 (.Z (n_580), .A (n_2524), .B (n_2482));
AOI22_X1 i_175 (.ZN (n_542), .A1 (n_476), .A2 (n_541), .B1 (n_540), .B2 (n_537));
XNOR2_X1 i_174 (.ZN (result[15]), .A (n_476), .B (n_541));
XOR2_X1 i_173 (.Z (n_541), .A (n_537), .B (n_540));
OAI21_X1 i_172 (.ZN (n_540), .A (n_539), .B1 (n_474), .B2 (n_538));
NAND2_X1 i_171 (.ZN (n_539), .A1 (n_474), .A2 (n_538));
AOI22_X1 i_170 (.ZN (n_538), .A1 (n_467), .A2 (n_454), .B1 (n_455), .B2 (n_466));
XNOR2_X1 i_169 (.ZN (n_537), .A (n_504), .B (n_536));
XOR2_X1 i_168 (.Z (n_536), .A (n_520), .B (n_535));
XOR2_X1 i_167 (.Z (n_535), .A (n_2415), .B (n_2414));
XOR2_X1 i_166 (.Z (n_520), .A (n_505), .B (n_519));
XNOR2_X1 i_165 (.ZN (n_519), .A (n_2110), .B (n_2119));
AOI22_X1 i_164 (.ZN (n_505), .A1 (n_465), .A2 (n_462), .B1 (n_463), .B2 (n_464));
XOR2_X1 i_163 (.Z (n_504), .A (n_501), .B (n_503));
AOI22_X1 i_162 (.ZN (n_503), .A1 (n_435), .A2 (n_453), .B1 (n_502), .B2 (n_434));
INV_X1 i_161 (.ZN (n_502), .A (n_413));
XOR2_X1 i_160 (.Z (n_501), .A (n_2484), .B (n_2483));
AOI21_X1 i_159 (.ZN (n_476), .A (n_469), .B1 (n_475), .B2 (n_471));
XNOR2_X1 i_158 (.ZN (result[14]), .A (n_472), .B (n_475));
AOI21_X1 i_157 (.ZN (n_475), .A (n_474), .B1 (n_407), .B2 (n_473));
NOR2_X1 i_156 (.ZN (n_474), .A1 (n_407), .A2 (n_473));
OAI22_X1 i_155 (.ZN (n_473), .A1 (n_355), .A2 (n_369), .B1 (n_367), .B2 (n_368));
NAND2_X1 i_154 (.ZN (n_472), .A1 (n_470), .A2 (n_471));
NAND2_X1 i_153 (.ZN (n_471), .A1 (n_411), .A2 (n_468));
INV_X1 i_152 (.ZN (n_470), .A (n_469));
NOR2_X1 i_151 (.ZN (n_469), .A1 (n_411), .A2 (n_468));
XOR2_X1 i_150 (.Z (n_468), .A (n_454), .B (n_467));
XOR2_X1 i_149 (.Z (n_467), .A (n_455), .B (n_466));
XOR2_X1 i_148 (.Z (n_466), .A (n_462), .B (n_465));
XOR2_X1 i_147 (.Z (n_465), .A (n_463), .B (n_464));
AOI22_X1 i_146 (.ZN (n_464), .A1 (n_402), .A2 (n_391), .B1 (n_401), .B2 (n_396));
AOI22_X1 i_145 (.ZN (n_463), .A1 (n_380), .A2 (n_386), .B1 (n_377), .B2 (n_379));
XOR2_X1 i_144 (.Z (n_462), .A (n_2424), .B (n_2418));
AOI22_X1 i_143 (.ZN (n_455), .A1 (n_404), .A2 (n_405), .B1 (n_387), .B2 (n_403));
XOR2_X1 i_142 (.Z (n_454), .A (n_435), .B (n_453));
XOR2_X1 i_141 (.Z (n_453), .A (n_2506), .B (n_2502));
XNOR2_X1 i_140 (.ZN (n_435), .A (n_413), .B (n_434));
XNOR2_X1 i_139 (.ZN (n_434), .A (n_2501), .B (n_2489));
NAND2_X1 i_138 (.ZN (n_16), .A1 (inputA[2]), .A2 (inputB[13]));
AOI22_X1 i_137 (.ZN (n_413), .A1 (n_365), .A2 (n_412), .B1 (n_357), .B2 (n_364));
INV_X1 i_136 (.ZN (n_412), .A (n_366));
OAI22_X1 i_135 (.ZN (n_411), .A1 (n_353), .A2 (n_409), .B1 (n_410), .B2 (n_370));
INV_X1 i_134 (.ZN (n_410), .A (n_408));
XNOR2_X1 i_133 (.ZN (result[13]), .A (n_353), .B (n_409));
XOR2_X1 i_132 (.Z (n_409), .A (n_370), .B (n_408));
OAI21_X1 i_131 (.ZN (n_408), .A (n_407), .B1 (n_371), .B2 (n_406));
NAND2_X1 i_130 (.ZN (n_407), .A1 (n_371), .A2 (n_406));
XOR2_X1 i_129 (.Z (n_406), .A (n_404), .B (n_405));
AOI22_X1 i_128 (.ZN (n_405), .A1 (n_306), .A2 (n_321), .B1 (n_2170), .B2 (n_320));
XOR2_X1 i_127 (.Z (n_404), .A (n_387), .B (n_403));
XOR2_X1 i_126 (.Z (n_403), .A (n_391), .B (n_402));
XOR2_X1 i_125 (.Z (n_402), .A (n_396), .B (n_401));
XNOR2_X1 i_124 (.ZN (n_401), .A (n_2137), .B (n_2136));
XOR2_X1 i_123 (.Z (n_396), .A (n_2122), .B (n_2121));
XOR2_X1 i_122 (.Z (n_391), .A (n_2430), .B (n_2429));
XOR2_X1 i_121 (.Z (n_387), .A (n_380), .B (n_386));
XOR2_X1 i_120 (.Z (n_386), .A (n_2131), .B (n_2130));
XOR2_X1 i_119 (.Z (n_380), .A (n_377), .B (n_379));
OAI21_X1 i_118 (.ZN (n_379), .A (n_2171), .B1 (n_378), .B2 (n_2174));
INV_X1 i_117 (.ZN (n_378), .A (n_2182));
XOR2_X1 i_116 (.Z (n_377), .A (n_374), .B (n_2421));
NOR2_X1 i_115 (.ZN (n_374), .A1 (n_2423), .A2 (n_2420));
INV_X1 i_114 (.ZN (n_371), .A (n_350));
XNOR2_X1 i_113 (.ZN (n_370), .A (n_355), .B (n_369));
XNOR2_X1 i_112 (.ZN (n_369), .A (n_367), .B (n_368));
AOI22_X1 i_111 (.ZN (n_368), .A1 (n_326), .A2 (n_342), .B1 (n_324), .B2 (n_325));
XOR2_X1 i_110 (.Z (n_367), .A (n_365), .B (n_366));
AOI22_X1 i_109 (.ZN (n_366), .A1 (n_337), .A2 (n_341), .B1 (n_332), .B2 (n_336));
XOR2_X1 i_108 (.Z (n_365), .A (n_357), .B (n_364));
XNOR2_X1 i_107 (.ZN (n_364), .A (n_2436), .B (n_2432));
AOI22_X1 i_106 (.ZN (n_357), .A1 (n_356), .A2 (n_2187), .B1 (n_2188), .B2 (n_2196));
INV_X1 i_105 (.ZN (n_356), .A (n_299));
AOI22_X1 i_104 (.ZN (n_355), .A1 (n_323), .A2 (n_343), .B1 (n_354), .B2 (n_322));
INV_X1 i_103 (.ZN (n_354), .A (n_298));
OAI21_X1 i_102 (.ZN (n_353), .A (n_345), .B1 (n_352), .B2 (n_351));
INV_X1 i_101 (.ZN (n_352), .A (n_346));
XOR2_X1 i_100 (.Z (result[12]), .A (n_347), .B (n_351));
OAI21_X1 i_99 (.ZN (n_351), .A (n_350), .B1 (n_348), .B2 (n_349));
NAND2_X1 i_98 (.ZN (n_350), .A1 (n_348), .A2 (n_349));
OAI21_X1 i_97 (.ZN (n_349), .A (n_288), .B1 (n_253), .B2 (n_289));
INV_X1 i_96 (.ZN (n_348), .A (n_293));
NAND2_X1 i_95 (.ZN (n_347), .A1 (n_345), .A2 (n_346));
OR2_X1 i_94 (.ZN (n_346), .A1 (n_296), .A2 (n_344));
NAND2_X1 i_93 (.ZN (n_345), .A1 (n_296), .A2 (n_344));
XNOR2_X1 i_92 (.ZN (n_344), .A (n_323), .B (n_343));
XOR2_X1 i_91 (.Z (n_343), .A (n_326), .B (n_342));
XOR2_X1 i_90 (.Z (n_342), .A (n_337), .B (n_341));
XNOR2_X1 i_89 (.ZN (n_341), .A (n_2451), .B (n_2441));
XOR2_X1 i_88 (.Z (n_337), .A (n_332), .B (n_336));
XNOR2_X1 i_87 (.ZN (n_336), .A (n_2422), .B (n_335));
NAND2_X1 i_86 (.ZN (n_335), .A1 (inputB[3]), .A2 (inputA[9]));
XOR2_X1 i_85 (.Z (n_332), .A (n_2439), .B (n_2140));
AOI22_X1 i_84 (.ZN (n_15), .A1 (inputB[4]), .A2 (inputA[8]), .B1 (inputB[5]), .B2 (inputA[7]));
XOR2_X1 i_83 (.Z (n_326), .A (n_324), .B (n_325));
AOI21_X1 i_82 (.ZN (n_325), .A (n_2249), .B1 (n_2248), .B2 (n_2247));
AOI22_X1 i_81 (.ZN (n_324), .A1 (n_2208), .A2 (n_2205), .B1 (n_2206), .B2 (n_2207));
XNOR2_X1 i_80 (.ZN (n_323), .A (n_298), .B (n_322));
XOR2_X1 i_79 (.Z (n_322), .A (n_306), .B (n_321));
XOR2_X1 i_78 (.Z (n_321), .A (n_2170), .B (n_320));
OAI21_X1 i_77 (.ZN (n_320), .A (n_2433), .B1 (n_2434), .B2 (n_2529));
AOI22_X1 i_76 (.ZN (n_14), .A1 (inputA[1]), .A2 (inputB[11]), .B1 (inputA[0]), .B2 (inputB[12]));
XOR2_X1 i_75 (.Z (n_306), .A (n_299), .B (n_2187));
AOI22_X1 i_74 (.ZN (n_299), .A1 (n_248), .A2 (n_249), .B1 (n_247), .B2 (n_245));
AOI22_X1 i_73 (.ZN (n_298), .A1 (n_251), .A2 (n_297), .B1 (n_244), .B2 (n_250));
INV_X1 i_72 (.ZN (n_297), .A (n_252));
AOI22_X1 i_71 (.ZN (n_296), .A1 (n_243), .A2 (n_295), .B1 (n_294), .B2 (n_290));
XNOR2_X1 i_70 (.ZN (result[11]), .A (n_243), .B (n_295));
XOR2_X1 i_69 (.Z (n_295), .A (n_290), .B (n_294));
OAI21_X1 i_68 (.ZN (n_294), .A (n_293), .B1 (n_291), .B2 (n_292));
NAND2_X1 i_67 (.ZN (n_293), .A1 (n_291), .A2 (n_292));
AOI22_X1 i_66 (.ZN (n_292), .A1 (n_2259), .A2 (n_235), .B1 (n_2260), .B2 (n_2286));
INV_X1 i_65 (.ZN (n_291), .A (n_2319));
XNOR2_X1 i_64 (.ZN (n_290), .A (n_253), .B (n_289));
OAI21_X1 i_63 (.ZN (n_289), .A (n_288), .B1 (n_2204), .B2 (n_2246));
NAND2_X1 i_62 (.ZN (n_288), .A1 (n_2246), .A2 (n_2204));
XNOR2_X1 i_61 (.ZN (n_253), .A (n_251), .B (n_252));
AOI22_X1 i_60 (.ZN (n_252), .A1 (n_234), .A2 (n_220), .B1 (n_229), .B2 (n_233));
XOR2_X1 i_59 (.Z (n_251), .A (n_244), .B (n_250));
XNOR2_X1 i_58 (.ZN (n_250), .A (n_248), .B (n_249));
OAI22_X1 i_57 (.ZN (n_249), .A1 (n_232), .A2 (n_2241), .B1 (n_2195), .B2 (n_231));
XOR2_X1 i_56 (.Z (n_248), .A (n_245), .B (n_247));
OAI33_X1 i_55 (.ZN (n_247), .A1 (n_2314), .A2 (n_690), .A3 (n_1349), .B1 (n_2186)
    , .B2 (n_1219), .B3 (n_864));
OAI22_X1 i_54 (.ZN (n_245), .A1 (n_2289), .A2 (n_2288), .B1 (n_2290), .B2 (n_2203));
AOI22_X1 i_53 (.ZN (n_244), .A1 (n_2291), .A2 (n_2287), .B1 (n_2292), .B2 (n_2312));
OAI22_X1 i_52 (.ZN (n_243), .A1 (n_199), .A2 (n_241), .B1 (n_242), .B2 (n_236));
INV_X1 i_51 (.ZN (n_242), .A (n_240));
XNOR2_X1 i_50 (.ZN (result[10]), .A (n_199), .B (n_241));
XOR2_X1 i_49 (.Z (n_241), .A (n_236), .B (n_240));
OAI21_X1 i_48 (.ZN (n_240), .A (n_2319), .B1 (n_2335), .B2 (n_2320));
XNOR2_X1 i_47 (.ZN (n_236), .A (n_2259), .B (n_235));
XOR2_X1 i_46 (.Z (n_235), .A (n_220), .B (n_234));
XOR2_X1 i_45 (.Z (n_234), .A (n_229), .B (n_233));
XNOR2_X1 i_44 (.ZN (n_233), .A (n_232), .B (n_2241));
XNOR2_X1 i_43 (.ZN (n_232), .A (n_2195), .B (n_231));
NAND2_X1 i_42 (.ZN (n_231), .A1 (inputA[0]), .A2 (inputB[10]));
XNOR2_X1 i_41 (.ZN (n_229), .A (n_2233), .B (n_2214));
AOI22_X1 i_40 (.ZN (n_220), .A1 (n_2327), .A2 (n_2325), .B1 (n_2329), .B2 (n_2328));
AOI22_X1 i_39 (.ZN (n_199), .A1 (n_163), .A2 (n_198), .B1 (n_166), .B2 (n_197));
XNOR2_X1 i_38 (.ZN (result[9]), .A (n_163), .B (n_198));
XOR2_X1 i_37 (.Z (n_198), .A (n_166), .B (n_197));
XOR2_X1 i_36 (.Z (n_197), .A (n_2331), .B (n_2321));
OAI21_X1 i_35 (.ZN (n_166), .A (n_2336), .B1 (n_2372), .B2 (n_2337));
OAI22_X1 i_34 (.ZN (n_163), .A1 (n_160), .A2 (n_162), .B1 (n_134), .B2 (n_159));
XNOR2_X1 i_33 (.ZN (result[8]), .A (n_160), .B (n_162));
AOI22_X1 i_32 (.ZN (n_162), .A1 (n_120), .A2 (n_161), .B1 (n_108), .B2 (n_119));
INV_X1 i_31 (.ZN (n_161), .A (n_121));
XNOR2_X1 i_30 (.ZN (n_160), .A (n_134), .B (n_159));
AOI21_X1 i_29 (.ZN (n_159), .A (n_2337), .B1 (n_2349), .B2 (n_2338));
XOR2_X1 i_28 (.Z (n_134), .A (n_2373), .B (n_2381));
XOR2_X1 i_27 (.Z (result[7]), .A (n_120), .B (n_121));
AOI22_X1 i_26 (.ZN (n_121), .A1 (n_94), .A2 (n_95), .B1 (n_90), .B2 (n_93));
XOR2_X1 i_25 (.Z (n_120), .A (n_108), .B (n_119));
XOR2_X1 i_24 (.Z (n_119), .A (n_2355), .B (n_2350));
OAI21_X1 i_23 (.ZN (n_108), .A (n_2373), .B1 (n_2374), .B2 (n_2380));
XNOR2_X1 i_22 (.ZN (result[6]), .A (n_94), .B (n_95));
OAI22_X1 i_21 (.ZN (n_95), .A1 (n_46), .A2 (n_65), .B1 (n_55), .B2 (n_64));
XOR2_X1 i_20 (.Z (n_94), .A (n_90), .B (n_93));
OAI21_X1 i_19 (.ZN (n_93), .A (n_2355), .B1 (n_2364), .B2 (n_2356));
XOR2_X1 i_18 (.Z (n_90), .A (n_2379), .B (n_2375));
XNOR2_X1 i_17 (.ZN (result[5]), .A (n_46), .B (n_65));
XNOR2_X1 i_16 (.ZN (n_65), .A (n_55), .B (n_64));
XOR2_X1 i_15 (.Z (n_64), .A (n_2359), .B (n_2357));
NAND2_X1 i_14 (.ZN (n_13), .A1 (inputB[0]), .A2 (inputA[5]));
AOI21_X1 i_13 (.ZN (n_55), .A (n_2364), .B1 (n_2366), .B2 (n_2365));
NAND2_X1 i_12 (.ZN (n_12), .A1 (inputA[1]), .A2 (inputB[4]));
AOI22_X1 i_11 (.ZN (n_46), .A1 (n_43), .A2 (n_45), .B1 (n_36), .B2 (n_42));
XNOR2_X1 i_10 (.ZN (result[4]), .A (n_43), .B (n_45));
AOI21_X1 i_9 (.ZN (n_45), .A (n_44), .B1 (n_73), .B2 (n_78));
INV_X1 i_8 (.ZN (n_44), .A (n_72));
XOR2_X1 i_7 (.Z (n_43), .A (n_36), .B (n_42));
XNOR2_X1 i_6 (.ZN (n_42), .A (n_2363), .B (n_2362));
AOI22_X1 i_5 (.ZN (n_11), .A1 (inputA[1]), .A2 (inputB[3]), .B1 (inputB[2]), .B2 (inputA[2]));
NOR2_X1 i_4 (.ZN (n_10), .A1 (n_61), .A2 (n_9));
NAND2_X1 i_3 (.ZN (n_9), .A1 (inputA[2]), .A2 (inputB[3]));
OAI21_X1 i_2 (.ZN (n_36), .A (n_2366), .B1 (n_2371), .B2 (n_2367));
NOR2_X1 i_1 (.ZN (result[1]), .A1 (n_51), .A2 (n_3));
AOI22_X1 i_0 (.ZN (n_3), .A1 (inputA[0]), .A2 (inputB[1]), .B1 (inputA[1]), .B2 (inputB[0]));

endmodule //datapath

module multiplyTimes (inputA, inputB, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;


datapath i_0 (.result ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32], result[31], 
    result[30], result[29], result[28], result[27], result[26], result[25], result[24], 
    result[23], result[22], result[21], result[20], result[19], result[18], result[17], 
    result[16], result[15], result[14], result[13], result[12], result[11], result[10], 
    result[9], result[8], result[7], result[6], result[5], result[4], result[3], 
    result[2], result[1], result[0]}), .inputA ({inputA[31], inputA[30], inputA[29], 
    inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], inputA[22], 
    inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], inputA[15], 
    inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], inputA[8], 
    inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], 
    inputA[0]}), .inputB ({inputB[31], inputB[30], inputB[29], inputB[28], inputB[27], 
    inputB[26], inputB[25], inputB[24], inputB[23], inputB[22], inputB[21], inputB[20], 
    inputB[19], inputB[18], inputB[17], inputB[16], inputB[15], inputB[14], inputB[13], 
    inputB[12], inputB[11], inputB[10], inputB[9], inputB[8], inputB[7], inputB[6], 
    inputB[5], inputB[4], inputB[3], inputB[2], inputB[1], inputB[0]}));

endmodule //multiplyTimes

module integrationMult (clk, reset, en, inputA, inputB, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n_tid1_3;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .en (en), .inp ({
    \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , 
    \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , 
    \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , 
    \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , 
    \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset), .clk_CTS_1_PP_0 (CTS_n_tid1_3));
registerNbits__2_8 outB (.out ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32]}), .clk_CTS_1_PP_0 (CTS_n_tid1_3)
    , .en (en), .inp ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , 
    \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , 
    \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , 
    \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , 
    \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , 
    \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , 
    \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTS_1_PP_1 (clk));
registerNbits__2_5 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTS_1_PP_0 (CTS_n_tid1_3));
registerNbits__2_2 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], 
    inputA[29], inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], 
    inputA[22], inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
    inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], 
    inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], 
    inputA[1], inputA[0]}), .reset (reset), .clk_CTS_1_PP_0 (CTS_n_tid1_3));
multiplyTimes mult (.result ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , 
    \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , 
    \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , 
    \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , 
    \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , 
    \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , 
    \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , 
    \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , 
    \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , 
    \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , 
    \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , 
    \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , 
    \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .inputA ({\A_reg[31] , \A_reg[30] , 
    \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , 
    \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , 
    \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , 
    \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , 
    \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] }), .inputB ({\B_reg[31] , 
    \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , \B_reg[25] , 
    \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , \B_reg[19] , 
    \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , \B_reg[13] , 
    \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , 
    \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }));

endmodule //integrationMult


