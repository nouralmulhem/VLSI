/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sun Dec 18 18:27:35 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 993135807 */

module fullAdder__1_185(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(cin), .A2(x), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(y), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(cin), .A2(x), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_3), .A2(y), .A3(n_0_0), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(y), .B1(n_0_3), .B2(n_0_0), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_182(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_179(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_176(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_173(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(y), .B(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
endmodule

module fullAdder__1_170(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   INV_X1 i_0_0 (.A(cin), .ZN(n_0_0));
   BUF_X1 i_0_1 (.A(n_0_2), .Z(n_0_1));
   INV_X1 i_0_2 (.A(n_0_7), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_3), .B1(n_0_4), .B2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_3));
   NOR2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(y), .ZN(n_0_5));
   OAI21_X1 i_0_7 (.A(n_0_6), .B1(x), .B2(n_0_9), .ZN(sum));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(n_0_0), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(n_0_1), .ZN(n_0_9));
endmodule

module fullAdder__1_167(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(x), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   XNOR2_X1 i_0_4 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_164(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_161(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_158(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_0), .B2(n_0_2), .ZN(cout));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(n_0_3), .ZN(sum));
   NAND2_X1 i_0_5 (.A1(n_0_6), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_7), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_155(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_152(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_149(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_146(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   XNOR2_X1 i_0_2 (.A(y), .B(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(x), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_3), .A2(x), .B1(n_0_4), .B2(n_0_1), .ZN(sum));
endmodule

module fullAdder__1_143(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_140(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_137(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_134(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_131(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_128(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_125(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_122(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_119(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_116(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_113(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_110(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_107(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_104(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_101(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_98(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_95(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_92(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_186(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_185 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_182 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_179 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_176 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_173 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_170 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_167 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_164 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_161 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_158 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_155 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_152 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_149 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_146 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_143 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_140 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_137 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_134 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_131 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_128 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_125 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_122 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_119 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_116 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_113 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_110 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_107 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_104 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_101 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_98 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(c1[2]));
   fullAdder__1_95 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(c1[1]));
   halfAdder__1_92 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_282(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NOR2_X1 i_0_2 (.A1(cin), .A2(x), .ZN(n_0_1));
   AND2_X1 i_0_3 (.A1(cin), .A2(x), .ZN(n_0_3));
   OR3_X1 i_0_5 (.A1(y), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   OAI21_X1 i_0_6 (.A(y), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_279(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_276(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_273(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_270(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_4), .B2(n_0_10), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_6), .A2(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_3), .A2(x), .A3(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(y), .ZN(n_0_5));
   OAI21_X1 i_0_8 (.A(n_0_10), .B1(n_0_7), .B2(n_0_9), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(y), .A2(cin), .ZN(n_0_8));
   NOR2_X1 i_0_11 (.A1(y), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(x), .ZN(n_0_10));
endmodule

module fullAdder__1_267(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_264(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_261(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_258(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_255(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(x), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   XNOR2_X1 i_0_4 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_252(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;

   INV_X1 i_0_0 (.A(x), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(cin), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_3), .ZN(cout));
   AOI21_X1 i_0_3 (.A(y), .B1(x), .B2(cin), .ZN(n_0_2));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(sum));
   NAND3_X1 i_0_6 (.A1(n_0_11), .A2(n_0_7), .A3(n_0_5), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(x), .A2(n_0_9), .A3(n_0_6), .ZN(n_0_5));
   OR2_X1 i_0_8 (.A1(y), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_10), .A2(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(n_0_9), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(x), .ZN(n_0_10));
   NAND2_X1 i_0_13 (.A1(n_0_0), .A2(n_0_12), .ZN(n_0_11));
   NOR2_X1 i_0_14 (.A1(y), .A2(n_0_13), .ZN(n_0_12));
   INV_X1 i_0_15 (.A(n_0_1), .ZN(n_0_13));
endmodule

module fullAdder__1_249(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_246(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_243(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_7), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(x), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(n_0_10), .B1(n_0_6), .B2(n_0_8), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(x), .A2(n_0_9), .ZN(n_0_7));
   NOR2_X1 i_0_10 (.A1(x), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_240(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_237(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_234(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_231(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_228(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_225(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_222(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_219(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_216(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_210(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_207(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_204(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_201(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_198(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_195(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_192(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_189(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_283(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_282 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_279 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_276 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_273 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_270 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_267 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_264 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_261 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_258 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_255 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_252 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_249 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_246 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_243 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_240 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_237 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_234 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_231 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_228 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_225 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_222 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_219 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_216 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_213 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_210 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_207 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_204 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_201 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_198 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_195 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_192 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_189 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_379(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_376(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_6), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(y), .A2(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_9), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_373(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_370(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_367(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_8), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_6), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_364(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_7), .B2(n_0_1), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(sum));
   AOI21_X1 i_0_4 (.A(x), .B1(n_0_6), .B2(n_0_5), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(x), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(y), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
endmodule

module fullAdder__1_361(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(cin), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_6), .ZN(sum));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(n_0_2), .ZN(n_0_8));
endmodule

module fullAdder__1_358(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   INV_X1 i_0_0 (.A(x), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_2));
   NOR2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   OAI21_X1 i_0_4 (.A(n_0_1), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_4), .A2(n_0_1), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(n_0_5), .ZN(n_0_6));
   AOI22_X1 i_0_8 (.A1(n_0_0), .A2(n_0_5), .B1(x), .B2(n_0_6), .ZN(sum));
endmodule

module fullAdder__1_355(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   OR2_X1 i_0_0 (.A1(y), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_1));
   AND3_X1 i_0_2 (.A1(x), .A2(n_0_0), .A3(n_0_1), .ZN(n_0_2));
   AOI21_X1 i_0_3 (.A(x), .B1(n_0_0), .B2(n_0_1), .ZN(n_0_3));
   NOR2_X1 i_0_4 (.A1(n_0_2), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_5 (.A(n_0_4), .B1(n_0_5), .B2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_352(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_349(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(x), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   XNOR2_X1 i_0_4 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_346(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(sum));
   AOI21_X1 i_0_3 (.A(x), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_5), .A2(x), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_7));
endmodule

module fullAdder__1_343(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_340(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_337(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_334(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_331(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_328(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_325(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_322(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_319(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_316(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_313(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_310(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_307(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_304(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_301(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_298(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_295(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_292(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_289(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_286(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_380(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_379 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_376 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_373 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_370 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_367 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_364 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_361 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_358 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_355 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_352 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_349 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_346 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_343 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_340 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_337 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_334 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_331 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_328 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_325 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_322 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_319 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_316 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_313 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_310 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_307 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_304 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_301 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_298 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_295 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_292 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_289 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_286 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_476(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(cin), .A2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(y), .A2(n_0_3), .ZN(n_0_2));
   OR2_X1 i_0_5 (.A1(cin), .A2(x), .ZN(n_0_3));
endmodule

module fullAdder__1_473(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_470(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_5), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_467(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;

   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(y), .A2(n_0_5), .A3(n_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_7), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_7));
   NAND2_X1 i_0_9 (.A1(n_0_9), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   NAND2_X1 i_0_12 (.A1(n_0_11), .A2(n_0_12), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
   INV_X1 i_0_14 (.A(cin), .ZN(n_0_12));
endmodule

module fullAdder__1_464(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_461(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_458(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_455(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(y), .B(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
endmodule

module fullAdder__1_452(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OR2_X1 i_0_0 (.A1(y), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND3_X1 i_0_2 (.A1(x), .A2(n_0_0), .A3(n_0_1), .ZN(n_0_2));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(x), .B1(n_0_0), .B2(n_0_1), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_449(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_446(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_443(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_440(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_437(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_434(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_431(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_428(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_425(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_422(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_419(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_416(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_413(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_410(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_407(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_404(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_401(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_398(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_395(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_392(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_389(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_386(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_383(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_477(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_476 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_473 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_470 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_467 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_464 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_461 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_458 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_455 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_452 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_449 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_446 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_443 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_440 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_437 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_434 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_431 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_428 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_425 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_422 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_419 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_416 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_413 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_410 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_407 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_404 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_401 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_398 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_395 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_392 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_389 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_386 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_383 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_573(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_570(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(y), .A2(n_0_3), .ZN(n_0_2));
   OR2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
endmodule

module fullAdder__1_567(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_6), .B1(n_0_2), .B2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   NAND3_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .A3(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_6), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_4), .B2(n_0_6), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_564(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_7), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(x), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(n_0_10), .B1(n_0_6), .B2(n_0_8), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(x), .A2(n_0_9), .ZN(n_0_7));
   NOR2_X1 i_0_10 (.A1(x), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_561(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_558(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_555(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_552(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_549(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_6), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
endmodule

module fullAdder__1_546(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_543(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_540(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_537(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_4), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_5), .ZN(sum));
   OAI21_X1 i_0_3 (.A(y), .B1(n_0_2), .B2(n_0_4), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(n_0_0), .B1(cin), .B2(x), .ZN(n_0_5));
endmodule

module fullAdder__1_534(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_531(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_528(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_525(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_522(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_519(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_516(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_513(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_510(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_507(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_504(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_501(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_498(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_495(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_492(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_489(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_486(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_483(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_480(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_574(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_573 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_570 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_567 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_564 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_561 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_558 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_555 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_552 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_549 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_546 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_543 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_540 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_537 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_534 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_531 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_528 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_525 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_522 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_519 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_516 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_513 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_510 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_507 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_504 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_501 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_498 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_495 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_492 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_489 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_486 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_483 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_480 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_670(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_667(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_664(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(y), .A2(n_0_3), .ZN(n_0_2));
   OR2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
endmodule

module fullAdder__1_661(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_7), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(y), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_7), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_8), .A2(n_0_7), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_5), .A2(n_0_6), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(x), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
endmodule

module fullAdder__1_658(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_655(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_6), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_652(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_649(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_646(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_643(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   INV_X1 i_0_0 (.A(x), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(cin), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_0), .A2(n_0_1), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(y), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_640(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_637(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_634(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_631(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_628(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   INV_X1 i_0_0 (.A(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_5), .ZN(cout));
   OAI21_X1 i_0_3 (.A(n_0_2), .B1(n_0_4), .B2(n_0_6), .ZN(sum));
   OAI21_X1 i_0_4 (.A(n_0_3), .B1(cin), .B2(x), .ZN(n_0_2));
   AOI21_X1 i_0_5 (.A(y), .B1(x), .B2(cin), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(n_0_0), .A2(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_625(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_622(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_619(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_616(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_613(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_610(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_607(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_604(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_601(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_598(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_595(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_592(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_589(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_586(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_583(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_580(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_577(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_671(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_670 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_667 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_664 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_661 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_658 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_655 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_652 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_649 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_646 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_643 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_640 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_637 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_634 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_631 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_628 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_625 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_622 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_619 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_616 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_613 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_610 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_607 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_604 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_601 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_598 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_595 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_592 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_589 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_586 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_583 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_580 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_577 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_767(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_764(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_761(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_758(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(y), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(x), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(cin), .ZN(n_0_5));
endmodule

module fullAdder__1_755(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_6), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_6), .A2(n_0_4), .A3(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_752(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_5), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_749(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_5), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_8), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_746(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_743(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_740(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_737(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(cin), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   NAND2_X1 i_0_8 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(n_0_7), .ZN(n_0_8));
   AOI22_X1 i_0_10 (.A1(n_0_6), .A2(n_0_8), .B1(x), .B2(n_0_7), .ZN(sum));
endmodule

module fullAdder__1_734(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(y), .B(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
endmodule

module fullAdder__1_731(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
   OAI22_X1 i_0_6 (.A1(n_0_3), .A2(cin), .B1(y), .B2(n_0_4), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(n_0_5), .ZN(n_0_6));
   AOI22_X1 i_0_8 (.A1(n_0_1), .A2(n_0_6), .B1(x), .B2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_728(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_725(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_722(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_719(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_716(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_713(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_710(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_707(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_704(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_701(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_698(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_695(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_692(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_689(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_686(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_683(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_680(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_677(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_674(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_768(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_767 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_764 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_761 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_758 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_755 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_752 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_749 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_746 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_743 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_740 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_737 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_734 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_731 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_728 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_725 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_722 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_719 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_716 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_713 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_710 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_707 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_704 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_701 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_698 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_695 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_692 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_689 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_686 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_683 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_680 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_677 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_674 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_864(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_861(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_858(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_855(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_852(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(n_0_1), .A2(y), .A3(n_0_2), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(n_0_7), .ZN(n_0_2));
   NAND3_X1 i_0_4 (.A1(n_0_8), .A2(n_0_5), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(cout));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   OAI21_X1 i_0_12 (.A(y), .B1(x), .B2(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_849(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_846(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_5), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_8), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_843(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_840(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_837(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_834(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_831(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_828(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(n_0_3), .B1(n_0_1), .B2(y), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(cin), .ZN(n_0_2));
   OR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_3));
   OR2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_5));
   AND3_X1 i_0_7 (.A1(n_0_4), .A2(x), .A3(n_0_5), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(x), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_7));
   NOR2_X1 i_0_9 (.A1(n_0_6), .A2(n_0_7), .ZN(sum));
endmodule

module fullAdder__1_825(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_822(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_819(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_816(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_813(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_810(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_807(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_804(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_801(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_798(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_795(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_792(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_789(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_786(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_783(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_780(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_777(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_774(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_771(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_865(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_864 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_861 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_858 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_855 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_852 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_849 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_846 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_843 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_840 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_837 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_834 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_831 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_828 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_825 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_822 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_819 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_816 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_813 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_810 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_807 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_804 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_801 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_798 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_795 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_792 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_789 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_786 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_783 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_780 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_777 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_774 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_771 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_961(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_958(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_955(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_952(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_949(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_946(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(n_0_1), .A2(y), .A3(n_0_5), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(x), .ZN(n_0_2));
   OAI21_X1 i_0_4 (.A(n_0_8), .B1(n_0_4), .B2(n_0_6), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_7), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_8));
   OAI21_X1 i_0_10 (.A(n_0_9), .B1(n_0_10), .B2(n_0_11), .ZN(cout));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   NOR2_X1 i_0_12 (.A1(x), .A2(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(y), .ZN(n_0_11));
endmodule

module fullAdder__1_943(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_940(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_8), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_937(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_934(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_931(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_928(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_2));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_3));
   OAI21_X1 i_0_4 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_5 (.A(x), .ZN(n_0_5));
   INV_X1 i_0_6 (.A(cin), .ZN(n_0_6));
   OAI21_X1 i_0_7 (.A(n_0_4), .B1(n_0_5), .B2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_8 (.A1(n_0_1), .A2(n_0_0), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(n_0_7), .ZN(n_0_8));
   AOI22_X1 i_0_10 (.A1(n_0_5), .A2(n_0_8), .B1(x), .B2(n_0_7), .ZN(sum));
endmodule

module fullAdder__1_925(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_922(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_919(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_916(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OR2_X1 i_0_0 (.A1(y), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND3_X1 i_0_2 (.A1(n_0_0), .A2(x), .A3(n_0_1), .ZN(n_0_2));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(x), .B1(n_0_0), .B2(n_0_1), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_913(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_910(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_907(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_904(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_901(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_898(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_895(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_892(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_889(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_886(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_883(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_880(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_877(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_874(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_871(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_868(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_962(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_961 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_958 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_955 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_952 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_949 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_946 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_943 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_940 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_937 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_934 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_931 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_928 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_925 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_922 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_919 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_916 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_913 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_910 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_907 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_904 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_901 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_898 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_895 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_892 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_889 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_886 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_883 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_880 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_877 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_874 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_871 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_868 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1058(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1055(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1052(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1049(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1046(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1043(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1040(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND3_X1 i_0_3 (.A1(x), .A2(n_0_5), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_1037(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1034(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1031(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1028(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1025(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   AOI21_X1 i_0_0 (.A(n_0_2), .B1(n_0_5), .B2(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(n_0_1), .ZN(n_0_0));
   OAI21_X1 i_0_3 (.A(n_0_5), .B1(n_0_3), .B2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(y), .ZN(n_0_5));
   OAI21_X1 i_0_8 (.A(y), .B1(n_0_8), .B2(n_0_7), .ZN(n_0_6));
   NOR2_X1 i_0_9 (.A1(x), .A2(n_0_10), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(n_0_9), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(x), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_1022(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_3 (.A(y), .B1(x), .B2(cin), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1019(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_3 (.A(y), .B1(x), .B2(cin), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1016(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_1013(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1010(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1007(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_0;
   wire n_0_1;
   wire n_0_3;
   wire n_0_5;
   wire n_0_2;
   wire n_0_9;
   wire n_0_4;

   AOI21_X1 i_0_0 (.A(n_0_2), .B1(n_0_8), .B2(n_0_4), .ZN(cout));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_1 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_0), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_4 (.A(y), .B1(x), .B2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_3));
   OAI21_X1 i_0_6 (.A(y), .B1(n_0_9), .B2(n_0_2), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_10 (.A(n_0_4), .ZN(n_0_9));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_4));
endmodule

module fullAdder__1_1004(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1001(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_998(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_995(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_992(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_989(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_986(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_983(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_980(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_977(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_974(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_971(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_968(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_965(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1059(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1058 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1055 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1052 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1049 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1046 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1043 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1040 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1037 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1034 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1031 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1028 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1025 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1022 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1019 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1016 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1013 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1010 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1007 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1004 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1001 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_998 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_995 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_992 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_989 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_986 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_983 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_980 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_977 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_974 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_971 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_968 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_965 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1155(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1152(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1149(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1146(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1143(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1140(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   AOI21_X1 i_0_0 (.A(n_0_2), .B1(n_0_5), .B2(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(n_0_1), .ZN(n_0_0));
   OAI21_X1 i_0_3 (.A(n_0_5), .B1(n_0_3), .B2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(y), .ZN(n_0_5));
   OAI21_X1 i_0_8 (.A(y), .B1(n_0_7), .B2(n_0_9), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(n_0_10), .ZN(n_0_8));
   NOR2_X1 i_0_11 (.A1(x), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_1137(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1134(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1131(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1128(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1125(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1122(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1119(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(n_0_1), .A2(y), .A3(n_0_2), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(n_0_7), .ZN(n_0_2));
   NAND3_X1 i_0_4 (.A1(n_0_8), .A2(n_0_5), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(cout));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   OAI21_X1 i_0_12 (.A(y), .B1(x), .B2(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_1116(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_1113(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NOR2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(y), .ZN(n_0_1));
   NAND2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_2));
   AOI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_0), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_0), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1110(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_6), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
endmodule

module fullAdder__1_1107(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1104(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1101(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1098(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1095(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1092(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1089(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1086(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1083(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1080(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1077(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1074(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1071(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1068(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1065(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1062(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1156(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1155 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1152 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1149 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1146 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1143 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1140 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1137 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1134 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1131 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1128 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1125 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1122 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1119 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1116 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1113 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1110 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1107 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1104 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1101 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1098 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1095 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1092 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1089 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1086 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1083 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1080 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1077 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1074 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1071 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1068 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1065 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1062 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1252(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1249(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1246(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1243(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1240(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1237(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1234(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_3), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_10), .A2(n_0_7), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1231(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1228(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1225(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1222(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1219(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1216(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1210(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_1207(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1204(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(x), .A2(n_0_7), .A3(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_10), .A2(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(y), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_9), .A2(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(x), .ZN(n_0_10));
endmodule

module fullAdder__1_1201(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_1198(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1195(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1192(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1189(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1186(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1183(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1180(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1177(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1174(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1171(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1168(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1165(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1162(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1159(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1253(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1252 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1249 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1246 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1243 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1240 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1237 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1234 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1231 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1228 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1225 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1222 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1219 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1216 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1213 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1210 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1207 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1204 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1201 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1198 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1195 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1192 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1189 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1186 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1183 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1180 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1177 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1174 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1171 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1168 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1165 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1162 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1159 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1349(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1346(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1343(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1340(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1337(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1334(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1331(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_6), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_6), .A2(n_0_4), .A3(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_1328(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1325(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1322(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_3));
   AND2_X1 i_0_5 (.A1(y), .A2(n_0_3), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(y), .A2(n_0_3), .ZN(n_0_5));
   NOR3_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .A3(x), .ZN(n_0_6));
   OR2_X1 i_0_8 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(n_0_6), .B1(n_0_7), .B2(x), .ZN(sum));
endmodule

module fullAdder__1_1319(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1316(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1313(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1310(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1307(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1304(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_4), .A2(x), .A3(n_0_9), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
   OAI21_X1 i_0_9 (.A(n_0_11), .B1(n_0_8), .B2(n_0_10), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(n_0_9), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(cin), .ZN(n_0_9));
   NOR2_X1 i_0_12 (.A1(y), .A2(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
endmodule

module fullAdder__1_1301(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_5), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(y), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(cin), .ZN(n_0_6));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(sum));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_1), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(x), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(n_0_1), .ZN(n_0_10));
endmodule

module fullAdder__1_1298(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1295(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OR2_X1 i_0_0 (.A1(y), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND3_X1 i_0_2 (.A1(x), .A2(n_0_0), .A3(n_0_1), .ZN(n_0_2));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(x), .B1(n_0_0), .B2(n_0_1), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_1292(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   OR2_X1 i_0_4 (.A1(y), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_4));
   AND3_X1 i_0_6 (.A1(x), .A2(n_0_3), .A3(n_0_4), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(x), .B1(n_0_3), .B2(n_0_4), .ZN(n_0_6));
   NOR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_6), .ZN(sum));
endmodule

module fullAdder__1_1289(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1286(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1283(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1280(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1277(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1274(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1271(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1268(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1265(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1262(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1259(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1256(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1350(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1349 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1346 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1343 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1340 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1337 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1334 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1331 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1328 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1325 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1322 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1319 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1316 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1313 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1310 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1307 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1304 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1301 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1298 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1295 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1292 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1289 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1286 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1283 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1280 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1277 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1274 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1271 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1268 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1265 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1262 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1259 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1256 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1446(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1443(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1440(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1437(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1434(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1431(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1428(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1425(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1422(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(y), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_8), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_9), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_10), .A2(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   NOR2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1419(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1416(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1413(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1410(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1407(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1404(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1401(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   AOI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_9), .B2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(sum));
   NAND3_X1 i_0_4 (.A1(y), .A2(n_0_7), .A3(n_0_5), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_9), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_5), .A2(n_0_7), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(x), .A2(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1398(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   AOI21_X1 i_0_0 (.A(n_0_6), .B1(n_0_4), .B2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_2 (.A1(n_0_1), .A2(n_0_4), .A3(n_0_8), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(x), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(y), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(y), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_1395(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND3_X1 i_0_8 (.A1(x), .A2(n_0_8), .A3(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(y), .A2(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1392(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1389(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1386(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1383(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1380(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1377(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1374(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1371(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1368(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1365(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1362(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1359(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1356(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1353(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1447(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1446 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1443 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1440 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1437 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1434 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1431 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1428 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1425 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1422 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1419 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1416 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1413 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1410 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1407 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1404 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1401 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1398 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1395 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1392 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1389 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1386 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1383 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1380 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1377 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1374 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1371 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1368 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1365 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1362 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1359 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1356 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1353 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1543(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1540(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1537(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1534(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1531(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1528(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1525(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1522(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1519(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1516(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1513(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1510(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_3), .ZN(cout));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum));
   AOI21_X1 i_0_2 (.A(x), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_4), .A2(x), .A3(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_1507(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1504(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1501(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_5), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1498(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1495(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_6), .B1(n_0_2), .B2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   NAND3_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .A3(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_6), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_4), .B2(n_0_6), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1492(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_5), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   OAI21_X1 i_0_3 (.A(n_0_2), .B1(n_0_4), .B2(n_0_6), .ZN(sum));
   OAI21_X1 i_0_4 (.A(n_0_3), .B1(cin), .B2(x), .ZN(n_0_2));
   AOI21_X1 i_0_5 (.A(y), .B1(x), .B2(cin), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(n_0_0), .A2(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_1489(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1486(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1483(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1480(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1477(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1474(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1471(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1468(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1465(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1462(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1459(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1456(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1453(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1450(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1544(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1543 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1540 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1537 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1534 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1531 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1528 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1525 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1522 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1519 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1516 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1513 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1510 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1507 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1504 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1501 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1498 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1495 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1492 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1489 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1486 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1483 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1480 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1477 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1474 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1471 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1468 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1465 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1462 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1459 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1456 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1453 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1450 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1640(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1637(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1634(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1631(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1628(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1625(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1622(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1619(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1616(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1613(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1610(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_5), .ZN(n_0_1));
   NAND3_X1 i_0_5 (.A1(n_0_4), .A2(n_0_9), .A3(n_0_7), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(x), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_1607(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1604(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1601(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   INV_X1 i_0_0 (.A(x), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(cin), .ZN(n_0_1));
   OAI21_X1 i_0_2 (.A(n_0_5), .B1(n_0_6), .B2(n_0_2), .ZN(cout));
   NOR2_X1 i_0_3 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_7), .ZN(sum));
   NAND3_X1 i_0_5 (.A1(n_0_4), .A2(n_0_6), .A3(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_0), .A2(n_0_1), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
   NAND3_X1 i_0_9 (.A1(n_0_8), .A2(y), .A3(n_0_9), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_0), .A2(cin), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(x), .A2(n_0_1), .ZN(n_0_9));
endmodule

module fullAdder__1_1598(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1595(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1592(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1589(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_8), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1586(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1583(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_3 (.A(y), .B1(x), .B2(cin), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1580(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   OR2_X1 i_0_3 (.A1(x), .A2(n_0_1), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_1), .ZN(n_0_4));
   NAND3_X1 i_0_6 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_5));
   AND2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_5), .B1(n_0_6), .B2(y), .ZN(sum));
endmodule

module fullAdder__1_1577(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1574(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1571(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1568(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1565(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1562(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1559(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1556(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1553(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1550(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1547(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1641(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1640 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1637 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1634 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1631 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1628 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1625 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1622 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1619 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1616 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1613 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1610 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1607 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1604 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1601 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1598 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1595 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1592 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1589 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1586 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1583 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1580 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1577 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1574 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1571 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1568 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1565 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1562 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1559 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1556 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1553 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1550 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1547 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1737(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1734(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1731(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1728(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1725(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1722(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1719(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1716(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1713(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1710(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1707(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1704(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1701(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1698(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1695(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1692(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(n_0_1), .A2(y), .A3(n_0_2), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(n_0_7), .ZN(n_0_2));
   NAND3_X1 i_0_4 (.A1(n_0_8), .A2(n_0_5), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(cout));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   OAI21_X1 i_0_12 (.A(y), .B1(x), .B2(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_1689(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   AOI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_9), .B2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(sum));
   NAND3_X1 i_0_4 (.A1(y), .A2(n_0_7), .A3(n_0_5), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_9), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_7), .A2(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1686(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1683(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1680(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1677(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_5;
   wire n_0_4;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_6;
   wire n_0_7;
   wire n_0_9;
   wire n_0_8;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;

   OAI21_X1 i_0_0 (.A(n_0_4), .B1(n_0_0), .B2(n_0_8), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_5), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_12), .A2(n_0_11), .ZN(n_0_5));
   NAND2_X1 i_0_3 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_4 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_7), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(n_0_12), .A2(n_0_6), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_9), .A2(n_0_10), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_8), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_12 (.A1(y), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(cin), .ZN(n_0_11));
   INV_X1 i_0_14 (.A(x), .ZN(n_0_12));
endmodule

module fullAdder__1_1674(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   AND2_X1 i_0_3 (.A1(x), .A2(n_0_1), .ZN(n_0_3));
   NOR2_X1 i_0_5 (.A1(x), .A2(n_0_1), .ZN(n_0_4));
   NOR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_4), .A3(y), .ZN(n_0_5));
   OR2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(n_0_5), .B1(y), .B2(n_0_6), .ZN(sum));
endmodule

module fullAdder__1_1671(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_6), .A2(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_6), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_11), .A2(n_0_9), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(x), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_10), .A2(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(y), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   NAND2_X1 i_0_12 (.A1(n_0_11), .A2(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(y), .ZN(n_0_11));
endmodule

module fullAdder__1_1668(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1665(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1662(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1659(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1656(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1653(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1650(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1647(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1644(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1738(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1737 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1734 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1731 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1728 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1725 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1722 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1719 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1716 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1713 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1710 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1707 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1704 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1701 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1698 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1695 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1692 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1689 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1686 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1683 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1680 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1677 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1674 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1671 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1668 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1665 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1662 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1659 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1656 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1653 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1650 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1647 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1644 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1834(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1831(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1828(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1825(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1822(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1819(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1816(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1813(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1810(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1807(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1804(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1801(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1798(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_7), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_8), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_6), .A2(n_0_10), .A3(n_0_9), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1795(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1792(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1789(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1786(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(y), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_10), .A2(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_11), .A2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_9), .A2(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(x), .A2(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(n_0_10), .A2(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(x), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(y), .ZN(n_0_11));
endmodule

module fullAdder__1_1783(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_5), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_8), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1780(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1777(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0_10), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND3_X1 i_0_8 (.A1(x), .A2(n_0_8), .A3(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(y), .A2(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1774(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_1771(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   OR2_X1 i_0_4 (.A1(y), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_4));
   AND3_X1 i_0_6 (.A1(x), .A2(n_0_3), .A3(n_0_4), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(x), .B1(n_0_3), .B2(n_0_4), .ZN(n_0_6));
   NOR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_6), .ZN(sum));
endmodule

module fullAdder__1_1768(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1765(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1762(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1759(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_11), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
endmodule

module fullAdder__1_1756(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_1753(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1750(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1747(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_1744(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1741(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1835(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1834 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1831 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1828 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1825 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1822 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1819 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1816 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1813 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1810 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1807 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1804 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1801 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1798 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1795 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1792 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1789 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1786 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1783 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1780 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1777 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1774 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1771 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1768 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1765 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1762 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1759 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1756 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1753 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1750 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1747 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1744 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1741 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_1931(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1928(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1925(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1922(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1919(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1916(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1913(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1910(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1907(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1904(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1901(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1898(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1895(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1892(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_7), .A3(n_0_5), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_9), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_7), .A2(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1889(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_10), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_9), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
   NAND2_X1 i_0_12 (.A1(y), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(cin), .ZN(n_0_11));
endmodule

module fullAdder__1_1886(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1883(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1880(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1877(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_5), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1874(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1871(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1868(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1865(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   OAI21_X1 i_0_0 (.A(n_0_8), .B1(n_0_0), .B2(n_0_10), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_9), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(n_0_1), .ZN(n_0_5));
   OAI21_X1 i_0_7 (.A(y), .B1(n_0_5), .B2(n_0_2), .ZN(n_0_6));
   NAND3_X1 i_0_8 (.A1(n_0_3), .A2(n_0_4), .A3(n_0_1), .ZN(n_0_7));
   NAND2_X1 i_0_9 (.A1(n_0_6), .A2(n_0_7), .ZN(sum));
   BUF_X1 i_0_10 (.A(n_0_1), .Z(n_0_8));
   BUF_X1 i_0_11 (.A(n_0_3), .Z(n_0_9));
   BUF_X1 i_0_12 (.A(n_0_4), .Z(n_0_10));
endmodule

module fullAdder__1_1862(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1859(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1856(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1853(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   OR2_X1 i_0_4 (.A1(y), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_4));
   AND3_X1 i_0_6 (.A1(x), .A2(n_0_3), .A3(n_0_4), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(x), .B1(n_0_3), .B2(n_0_4), .ZN(n_0_6));
   NOR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_6), .ZN(sum));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(y), .ZN(n_0_2));
endmodule

module fullAdder__1_1850(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1847(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1844(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   XNOR2_X1 i_0_8 (.A(y), .B(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_1841(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_1838(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_1932(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_1931 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_1928 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_1925 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_1922 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_1919 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_1916 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_1913 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_1910 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_1907 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_1904 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1901 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1898 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1895 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1892 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1889 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1886 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1883 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1880 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1877 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1874 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1871 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1868 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1865 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1862 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1859 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1856 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1853 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1850 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1847 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1844 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1841 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1838 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2028(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2025(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2022(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2019(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2016(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2013(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2010(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2007(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2004(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2001(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1998(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1995(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1992(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1989(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1986(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1983(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1980(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_1977(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1974(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1971(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1968(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1965(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_6), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_8), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_6), .A2(n_0_9), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_1962(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1959(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND3_X1 i_0_8 (.A1(x), .A2(n_0_8), .A3(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(y), .A2(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_1956(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1953(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   OAI21_X1 i_0_4 (.A(y), .B1(x), .B2(cin), .ZN(n_0_2));
endmodule

module fullAdder__1_1950(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1947(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1944(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_1941(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_6), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_6), .A2(n_0_4), .A3(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_1938(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module halfAdder__1_1935(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2029(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2028 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2025 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2022 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2019 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2016 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2013 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2010 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2007 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2004 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2001 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_1998 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_1995 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_1992 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_1989 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_1986 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_1983 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_1980 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_1977 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_1974 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_1971 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_1968 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_1965 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_1962 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_1959 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_1956 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_1953 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_1950 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_1947 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_1944 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_1941 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_1938 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_1935 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2125(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2122(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2119(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2116(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2113(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2110(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2107(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2104(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2101(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2098(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2095(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2092(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2089(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2086(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2083(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2080(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2077(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2074(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2071(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2068(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2065(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND3_X1 i_0_1 (.A1(n_0_1), .A2(y), .A3(n_0_2), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(n_0_7), .ZN(n_0_2));
   NAND3_X1 i_0_4 (.A1(n_0_5), .A2(n_0_8), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(cout));
   NAND2_X1 i_0_11 (.A1(x), .A2(cin), .ZN(n_0_9));
   OAI21_X1 i_0_12 (.A(y), .B1(x), .B2(cin), .ZN(n_0_10));
endmodule

module fullAdder__1_2062(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2059(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND3_X1 i_0_3 (.A1(x), .A2(n_0_5), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_8), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_7), .A2(n_0_6), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(y), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
endmodule

module fullAdder__1_2056(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2053(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   AOI21_X1 i_0_0 (.A(n_0_2), .B1(n_0_8), .B2(n_0_4), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_4), .ZN(n_0_1));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_5), .A2(n_0_8), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
endmodule

module fullAdder__1_2050(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2047(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2044(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_2041(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2038(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2035(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_2032(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2126(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2125 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2122 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2119 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2116 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2113 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2110 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2107 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2104 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2101 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2098 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2095 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2092 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2089 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2086 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2083 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2080 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2077 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2074 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2071 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2068 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2065 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2062 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2059 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2056 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2053 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2050 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2047 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2044 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2041 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2038 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2035 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2032 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2222(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2219(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2216(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2210(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2207(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2204(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2201(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2198(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2195(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2192(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2189(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2186(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2183(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2180(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2177(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2174(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2171(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2168(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2165(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2162(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2159(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2156(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_6), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_6), .A2(n_0_4), .A3(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(y), .ZN(n_0_6));
endmodule

module fullAdder__1_2153(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2150(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2147(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2144(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2141(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_11), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
endmodule

module fullAdder__1_2138(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2135(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2132(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   AND2_X1 i_0_3 (.A1(y), .A2(n_0_1), .ZN(n_0_3));
   NOR2_X1 i_0_5 (.A1(y), .A2(n_0_1), .ZN(n_0_4));
   NOR3_X1 i_0_6 (.A1(n_0_3), .A2(x), .A3(n_0_4), .ZN(n_0_5));
   OR2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(n_0_5), .B1(n_0_6), .B2(x), .ZN(sum));
endmodule

module halfAdder__1_2129(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2223(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2222 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2219 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2216 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2213 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2210 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2207 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2204 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2201 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2198 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2195 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2192 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2189 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2186 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2183 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2180 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2177 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2174 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2171 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2168 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2165 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2162 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2159 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2156 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2153 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2150 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2147 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2144 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2141 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2138 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2135 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2132 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2129 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2319(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2316(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2313(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2310(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2307(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2304(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2301(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2298(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2295(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2292(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2289(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2286(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2283(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2280(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2277(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2274(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2271(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2268(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2265(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2262(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2259(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2256(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2253(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2250(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2247(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_5), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(n_0_6), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(y), .A2(n_0_2), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_8), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_9), .A2(n_0_6), .A3(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(x), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(x), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2244(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(n_0_1), .A2(x), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2241(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   AOI21_X1 i_0_0 (.A(n_0_6), .B1(n_0_4), .B2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_5), .ZN(sum));
   NAND3_X1 i_0_2 (.A1(n_0_4), .A2(n_0_8), .A3(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(x), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(y), .ZN(n_0_4));
   OAI21_X1 i_0_7 (.A(y), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_2238(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2235(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2232(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2229(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_2226(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2320(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2319 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2316 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2313 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2310 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2307 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2304 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2301 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2298 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2295 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2292 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2289 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2286 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2283 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2280 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2277 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2274 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2271 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2268 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2265 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2262 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2259 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2256 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2253 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2250 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2247 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2244 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2241 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2238 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2235 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2232 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2229 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2226 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2416(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2413(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2410(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2407(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2404(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2401(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2398(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2395(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2392(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2389(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2386(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2383(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2380(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2377(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2374(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2371(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2368(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2365(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2362(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2359(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2356(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2353(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2350(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2347(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_10), .A2(n_0_7), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2344(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2341(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2338(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2335(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2332(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_2329(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2326(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_2323(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2417(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2416 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2413 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2410 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2407 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2404 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2401 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2398 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2395 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2392 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2389 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2386 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2383 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2380 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2377 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2374 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2371 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2368 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2365 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2362 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2359 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2356 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2353 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2350 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2347 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2344 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2341 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2338 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2335 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2332 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2329 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2326 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2323 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2513(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2510(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2507(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2504(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2501(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2498(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2495(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2492(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2489(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2486(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2483(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2480(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2477(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2474(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2471(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2468(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2465(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2462(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2459(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2456(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2453(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2450(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2447(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2444(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2441(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2438(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2435(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_8), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(y), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_2), .A2(y), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_7), .ZN(n_0_3));
   NAND3_X1 i_0_6 (.A1(n_0_5), .A2(n_0_9), .A3(n_0_8), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_7), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(x), .A2(cin), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(y), .ZN(n_0_9));
endmodule

module fullAdder__1_2432(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2429(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   OAI21_X1 i_0_4 (.A(y), .B1(x), .B2(cin), .ZN(n_0_2));
endmodule

module fullAdder__1_2426(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(y), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_0), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_1), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_1), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2423(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_2420(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2514(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2513 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2510 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2507 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2504 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2501 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2498 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2495 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2492 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2489 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2486 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2483 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2480 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2477 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2474 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2471 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2468 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2465 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2462 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2459 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2456 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2453 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2450 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2447 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2444 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2441 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2438 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2435 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2432 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2429 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2426 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2423 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2420 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2610(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2607(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2604(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2601(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2598(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2595(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2592(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2589(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2586(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2583(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2580(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2577(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2574(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2571(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2568(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2565(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2562(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2559(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2556(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2553(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2550(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2547(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2544(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2541(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2538(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2535(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2532(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module fullAdder__1_2529(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2526(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   OAI21_X1 i_0_0 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(x), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_2));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   AND2_X1 i_0_4 (.A1(y), .A2(n_0_2), .ZN(n_0_3));
   NOR2_X1 i_0_5 (.A1(y), .A2(n_0_2), .ZN(n_0_4));
   NOR3_X1 i_0_6 (.A1(n_0_3), .A2(x), .A3(n_0_4), .ZN(n_0_5));
   OR2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(n_0_5), .B1(n_0_6), .B2(x), .ZN(sum));
endmodule

module fullAdder__1_2523(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2520(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;

   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(x), .A2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(y), .ZN(n_0_3));
endmodule

module halfAdder__1_2517(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2611(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2610 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2607 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2604 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2601 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2598 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2595 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2592 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2589 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2586 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2583 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2580 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2577 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2574 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2571 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2568 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2565 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2562 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2559 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2556 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2553 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2550 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2547 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2544 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2541 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2538 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2535 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2532 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2529 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2526 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2523 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2520 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2517 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2707(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2704(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2701(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2698(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2695(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2692(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2689(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2686(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2683(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2680(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2677(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2674(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2671(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2668(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2665(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2662(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2659(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2656(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2653(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2650(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2647(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2644(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2641(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2638(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2635(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2632(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2629(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_7), .ZN(n_0_1));
   OAI21_X1 i_0_5 (.A(n_0_6), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(y), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_11), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
   NAND3_X1 i_0_9 (.A1(n_0_8), .A2(x), .A3(n_0_11), .ZN(n_0_7));
   NAND2_X1 i_0_10 (.A1(n_0_10), .A2(n_0_9), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
   NAND2_X1 i_0_13 (.A1(y), .A2(cin), .ZN(n_0_11));
endmodule

module fullAdder__1_2626(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2623(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2620(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NOR2_X1 i_0_0 (.A1(x), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(y), .ZN(n_0_1));
   NAND2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_2));
   AOI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_0_2), .ZN(cout));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_3), .B2(n_0_0), .ZN(n_0_4));
   OR3_X1 i_0_6 (.A1(n_0_3), .A2(n_0_0), .A3(y), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module fullAdder__1_2617(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder__1_2614(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2708(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2707 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2704 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2701 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2698 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2695 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2692 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2689 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2686 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2683 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2680 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2677 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2674 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2671 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2668 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2665 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2662 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2659 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2656 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2653 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2650 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2647 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2644 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2641 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2638 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2635 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2632 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2629 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2626 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2623 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2620 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2617 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2614 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2804(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2801(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2798(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2795(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2792(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2789(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2786(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2783(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2780(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2777(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2774(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2771(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2768(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2765(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2762(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2759(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2756(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2753(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2750(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2747(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2744(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2741(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2738(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_2735(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_6), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_11), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_9), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
endmodule

module fullAdder__1_2732(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2729(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2726(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2723(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   NAND2_X1 i_0_2 (.A1(n_0_5), .A2(n_0_1), .ZN(sum));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_8), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(x), .A2(n_0_9), .ZN(n_0_4));
   NAND3_X1 i_0_7 (.A1(n_0_7), .A2(n_0_10), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(x), .ZN(n_0_8));
   INV_X1 i_0_11 (.A(cin), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(y), .ZN(n_0_10));
endmodule

module fullAdder__1_2720(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(y), .ZN(n_0_0));
   OR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(x), .A2(cin), .ZN(n_0_2));
   OR2_X1 i_0_4 (.A1(y), .A2(cin), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y), .A2(cin), .ZN(n_0_4));
   AND3_X1 i_0_6 (.A1(x), .A2(n_0_3), .A3(n_0_4), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(x), .B1(n_0_3), .B2(n_0_4), .ZN(n_0_6));
   NOR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_6), .ZN(sum));
endmodule

module fullAdder__1_2717(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_2714(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   OR2_X1 i_0_2 (.A1(y), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(y), .A2(cin), .ZN(n_0_3));
   AND3_X1 i_0_5 (.A1(x), .A2(n_0_1), .A3(n_0_3), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_1), .B2(n_0_3), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_5), .ZN(sum));
endmodule

module halfAdder__1_2711(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__1_2805(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2804 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_2801 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_2798 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_2795 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_2792 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_2789 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_2786 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_2783 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_2780 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_2777 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_2774 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_2771 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_2768 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_2765 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_2762 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_2759 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_2756 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_2753 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_2750 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_2747 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_2744 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_2741 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_2738 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_2735 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(
      c1[8]));
   fullAdder__1_2732 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(
      c1[7]));
   fullAdder__1_2729 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(
      c1[6]));
   fullAdder__1_2726 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(
      c1[5]));
   fullAdder__1_2723 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(
      c1[4]));
   fullAdder__1_2720 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(
      c1[3]));
   fullAdder__1_2717 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(
      c1[2]));
   fullAdder__1_2714 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(
      c1[1]));
   halfAdder__1_2711 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module fullAdder__1_2(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_5(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_8(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_11(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_14(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_17(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_20(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_23(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_26(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_29(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_32(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_35(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_38(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_41(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_44(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_47(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_50(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_53(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_56(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_59(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_62(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_65(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__1_68(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   XNOR2_X1 i_0_3 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_1), .A2(n_0_3), .B1(x), .B2(n_0_4), .ZN(sum));
endmodule

module fullAdder__1_71(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_1));
   OAI21_X1 i_0_5 (.A(x), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(y), .A2(n_0_10), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_9), .ZN(n_0_5));
   NAND3_X1 i_0_8 (.A1(n_0_11), .A2(n_0_9), .A3(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_8), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(y), .A2(n_0_10), .ZN(n_0_9));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(x), .ZN(n_0_11));
endmodule

module fullAdder__1_74(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_5), .ZN(n_0_2));
   XNOR2_X1 i_0_4 (.A(y), .B(cin), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(x), .ZN(n_0_4));
   AOI22_X1 i_0_6 (.A1(n_0_4), .A2(n_0_3), .B1(x), .B2(n_0_2), .ZN(sum));
   BUF_X1 i_0_7 (.A(n_0_3), .Z(n_0_5));
endmodule

module fullAdder__1_77(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(x), .B2(cin), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(x), .A2(cin), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(sum));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_6), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_7), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(x), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(n_0_7), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y), .B(n_0_8), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(cin), .ZN(n_0_8));
endmodule

module fullAdder__1_80(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(y), .B(cin), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(x), .ZN(n_0_6));
endmodule

module fullAdder__1_83(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_4), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(sum));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_3 (.A(y), .B1(x), .B2(cin), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(n_0_2));
   OAI21_X1 i_0_5 (.A(y), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(x), .A2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module fullAdder__1_86(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   OR2_X1 i_0_3 (.A1(x), .A2(n_0_1), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(x), .A2(n_0_1), .ZN(n_0_4));
   NAND3_X1 i_0_6 (.A1(n_0_3), .A2(y), .A3(n_0_4), .ZN(n_0_5));
   AND2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_5), .B1(n_0_6), .B2(y), .ZN(sum));
endmodule

module fullAdder__1_89(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   AOI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_7), .B2(n_0_1), .ZN(cout));
   AOI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(x), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_4), .ZN(sum));
   INV_X1 i_0_4 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_6), .A2(x), .A3(n_0_5), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(x), .B1(n_0_6), .B2(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(y), .A2(cin), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(y), .ZN(n_0_8));
endmodule

module fullAdder__0_46(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_4), .A2(n_0_6), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_0), .A2(n_0_3), .ZN(sum));
   OAI21_X1 i_0_2 (.A(y), .B1(n_0_1), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   AOI21_X1 i_0_6 (.A(y), .B1(x), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_8 (.A1(x), .A2(cin), .ZN(n_0_6));
endmodule

module halfAdder__0_43(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder__0_47(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__1_2 fa31 (.x(a[32]), .y(b[31]), .cin(c[30]), .sum(s1[31]), 
      .cout(c1[31]));
   fullAdder__1_5 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__1_8 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__1_11 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__1_14 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__1_17 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__1_20 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__1_23 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__1_26 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__1_29 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__1_32 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__1_35 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__1_38 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__1_41 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__1_44 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__1_47 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__1_50 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__1_53 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__1_56 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__1_59 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__1_62 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__1_65 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__1_68 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__1_71 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(c1[8]));
   fullAdder__1_74 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(c1[7]));
   fullAdder__1_77 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(c1[6]));
   fullAdder__1_80 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(c1[5]));
   fullAdder__1_83 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(c1[4]));
   fullAdder__1_86 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(c1[3]));
   fullAdder__1_89 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(c1[2]));
   fullAdder__0_46 fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(c1[1]));
   halfAdder__0_43 ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module datapath(b, a, p_0);
   input [31:0]b;
   input [31:0]a;
   output [32:0]p_0;

   XOR2_X1 i_0 (.A(n_0), .B(n_193), .Z(p_0[6]));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_2), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_88), .B(n_124), .Z(p_0[12]));
   INV_X1 i_3 (.A(n_4), .ZN(p_0[13]));
   XOR2_X1 i_4 (.A(n_5), .B(n_9), .Z(n_4));
   NAND2_X1 i_5 (.A1(n_111), .A2(n_117), .ZN(n_5));
   XOR2_X1 i_6 (.A(n_6), .B(n_8), .Z(p_0[14]));
   NAND2_X1 i_7 (.A1(n_113), .A2(n_110), .ZN(n_6));
   XNOR2_X1 i_8 (.A(n_7), .B(n_11), .ZN(p_0[15]));
   AOI21_X1 i_9 (.A(n_112), .B1(n_8), .B2(n_110), .ZN(n_7));
   OAI21_X1 i_10 (.A(n_111), .B1(n_9), .B2(n_10), .ZN(n_8));
   OAI21_X1 i_11 (.A(n_89), .B1(n_124), .B2(n_90), .ZN(n_9));
   INV_X1 i_12 (.A(n_117), .ZN(n_10));
   NAND2_X1 i_13 (.A1(n_116), .A2(n_109), .ZN(n_11));
   INV_X1 i_14 (.A(n_12), .ZN(p_0[16]));
   XOR2_X1 i_15 (.A(n_13), .B(n_130), .Z(n_12));
   NAND2_X1 i_16 (.A1(n_20), .A2(n_107), .ZN(n_13));
   XOR2_X1 i_17 (.A(n_14), .B(n_18), .Z(p_0[17]));
   NAND2_X1 i_18 (.A1(n_106), .A2(n_108), .ZN(n_14));
   XNOR2_X1 i_19 (.A(n_17), .B(n_91), .ZN(p_0[18]));
   XNOR2_X1 i_20 (.A(n_16), .B(n_94), .ZN(p_0[19]));
   OAI21_X1 i_21 (.A(n_93), .B1(n_17), .B2(n_21), .ZN(n_16));
   AOI21_X1 i_22 (.A(n_105), .B1(n_18), .B2(n_108), .ZN(n_17));
   AOI21_X1 i_23 (.A(n_19), .B1(n_130), .B2(n_20), .ZN(n_18));
   INV_X1 i_24 (.A(n_107), .ZN(n_19));
   NAND2_X1 i_25 (.A1(n_132), .A2(n_131), .ZN(n_20));
   INV_X1 i_26 (.A(n_92), .ZN(n_21));
   XOR2_X1 i_27 (.A(n_101), .B(n_137), .Z(p_0[20]));
   INV_X1 i_28 (.A(n_26), .ZN(p_0[21]));
   XOR2_X1 i_29 (.A(n_27), .B(n_28), .Z(n_26));
   NAND2_X1 i_30 (.A1(n_139), .A2(n_104), .ZN(n_27));
   OAI21_X1 i_31 (.A(n_102), .B1(n_137), .B2(n_103), .ZN(n_28));
   XNOR2_X1 i_32 (.A(n_42), .B(n_41), .ZN(p_0[25]));
   NAND2_X1 i_33 (.A1(n_164), .A2(n_166), .ZN(n_41));
   NAND2_X1 i_34 (.A1(n_165), .A2(n_160), .ZN(n_42));
   INV_X1 i_35 (.A(n_64), .ZN(p_0[28]));
   XOR2_X1 i_36 (.A(n_65), .B(n_100), .Z(n_64));
   NAND2_X1 i_37 (.A1(n_99), .A2(n_192), .ZN(n_65));
   XNOR2_X1 i_38 (.A(n_67), .B(n_66), .ZN(p_0[29]));
   NAND2_X1 i_39 (.A1(n_182), .A2(n_181), .ZN(n_66));
   NAND2_X1 i_40 (.A1(n_98), .A2(n_192), .ZN(n_67));
   NAND2_X1 i_41 (.A1(n_69), .A2(n_68), .ZN(p_0[30]));
   NAND3_X1 i_42 (.A1(n_71), .A2(n_182), .A3(n_73), .ZN(n_68));
   NAND2_X1 i_43 (.A1(n_70), .A2(n_72), .ZN(n_69));
   NAND2_X1 i_44 (.A1(n_71), .A2(n_182), .ZN(n_70));
   NAND3_X1 i_45 (.A1(n_98), .A2(n_192), .A3(n_181), .ZN(n_71));
   INV_X1 i_46 (.A(n_73), .ZN(n_72));
   NAND2_X1 i_47 (.A1(n_204), .A2(n_180), .ZN(n_73));
   NAND2_X1 i_48 (.A1(n_74), .A2(n_77), .ZN(p_0[31]));
   NAND2_X1 i_49 (.A1(n_75), .A2(n_76), .ZN(n_74));
   NAND2_X1 i_50 (.A1(n_79), .A2(n_78), .ZN(n_75));
   INV_X1 i_51 (.A(n_82), .ZN(n_76));
   NAND3_X1 i_52 (.A1(n_79), .A2(n_82), .A3(n_78), .ZN(n_77));
   AOI21_X1 i_53 (.A(n_207), .B1(n_183), .B2(n_180), .ZN(n_78));
   NAND3_X1 i_54 (.A1(n_98), .A2(n_192), .A3(n_179), .ZN(n_79));
   NAND2_X1 i_55 (.A1(n_208), .A2(n_211), .ZN(n_82));
   OAI21_X1 i_56 (.A(n_189), .B1(n_98), .B2(n_203), .ZN(p_0[32]));
   NAND2_X1 i_57 (.A1(n_100), .A2(n_99), .ZN(n_98));
   OR2_X1 i_58 (.A1(a[28]), .A2(b[28]), .ZN(n_99));
   OAI21_X1 i_59 (.A(n_184), .B1(n_137), .B2(n_114), .ZN(n_100));
   NAND2_X1 i_60 (.A1(n_154), .A2(n_187), .ZN(n_114));
   NAND2_X1 i_61 (.A1(b[0]), .A2(a[0]), .ZN(n_15));
   NAND2_X1 i_62 (.A1(b[1]), .A2(a[1]), .ZN(n_22));
   NAND2_X1 i_63 (.A1(n_39), .A2(n_38), .ZN(n_193));
   XOR2_X1 i_217 (.A(b[0]), .B(a[0]), .Z(p_0[0]));
   NAND2_X1 i_64 (.A1(n_51), .A2(n_22), .ZN(n_194));
   XOR2_X1 i_65 (.A(n_194), .B(n_15), .Z(p_0[1]));
   NAND2_X1 i_66 (.A1(n_53), .A2(n_51), .ZN(n_195));
   NAND2_X1 i_67 (.A1(n_52), .A2(n_48), .ZN(n_196));
   XOR2_X1 i_68 (.A(n_195), .B(n_196), .Z(p_0[2]));
   NAND2_X1 i_69 (.A1(n_50), .A2(n_48), .ZN(n_197));
   NAND2_X1 i_70 (.A1(n_45), .A2(n_49), .ZN(n_198));
   XNOR2_X1 i_71 (.A(n_197), .B(n_198), .ZN(p_0[3]));
   NAND2_X1 i_72 (.A1(n_47), .A2(n_45), .ZN(n_199));
   NAND2_X1 i_73 (.A1(n_46), .A2(n_40), .ZN(n_200));
   XOR2_X1 i_74 (.A(n_199), .B(n_200), .Z(p_0[4]));
   NAND2_X1 i_75 (.A1(n_44), .A2(n_40), .ZN(n_201));
   NAND2_X1 i_76 (.A1(n_38), .A2(n_43), .ZN(n_202));
   XNOR2_X1 i_77 (.A(n_201), .B(n_202), .ZN(p_0[5]));
   NAND3_X1 i_78 (.A1(n_39), .A2(n_38), .A3(n_37), .ZN(n_205));
   NAND2_X1 i_79 (.A1(n_205), .A2(n_33), .ZN(n_206));
   NAND2_X1 i_80 (.A1(n_35), .A2(n_34), .ZN(n_210));
   XNOR2_X1 i_81 (.A(n_206), .B(n_210), .ZN(p_0[7]));
   NAND2_X1 i_82 (.A1(n_25), .A2(n_30), .ZN(n_1));
   XNOR2_X1 i_83 (.A(n_31), .B(n_1), .ZN(p_0[8]));
   BUF_X1 i_84 (.A(n_33), .Z(n_2));
   BUF_X1 i_85 (.A(n_37), .Z(n_3));
   XNOR2_X1 i_86 (.A(n_24), .B(n_23), .ZN(p_0[9]));
   NAND2_X1 i_87 (.A1(n_55), .A2(n_54), .ZN(n_23));
   NAND2_X1 i_88 (.A1(n_29), .A2(n_25), .ZN(n_24));
   NAND2_X1 i_89 (.A1(b[8]), .A2(a[8]), .ZN(n_25));
   NAND2_X1 i_90 (.A1(n_31), .A2(n_30), .ZN(n_29));
   NAND2_X1 i_91 (.A1(n_58), .A2(n_57), .ZN(n_30));
   OAI221_X1 i_92 (.A(n_34), .B1(n_36), .B2(n_33), .C1(n_36), .C2(n_32), 
      .ZN(n_31));
   NAND3_X1 i_93 (.A1(n_39), .A2(n_38), .A3(n_37), .ZN(n_32));
   NAND2_X1 i_94 (.A1(b[6]), .A2(a[6]), .ZN(n_33));
   NAND2_X1 i_95 (.A1(b[7]), .A2(a[7]), .ZN(n_34));
   INV_X1 i_96 (.A(n_36), .ZN(n_35));
   NOR2_X1 i_97 (.A1(b[7]), .A2(a[7]), .ZN(n_36));
   OR2_X1 i_98 (.A1(b[6]), .A2(a[6]), .ZN(n_37));
   OR2_X1 i_99 (.A1(b[5]), .A2(a[5]), .ZN(n_38));
   NAND3_X1 i_100 (.A1(n_44), .A2(n_43), .A3(n_40), .ZN(n_39));
   NAND2_X1 i_101 (.A1(b[4]), .A2(a[4]), .ZN(n_40));
   NAND2_X1 i_102 (.A1(b[5]), .A2(a[5]), .ZN(n_43));
   NAND3_X1 i_103 (.A1(n_47), .A2(n_46), .A3(n_45), .ZN(n_44));
   OR2_X1 i_104 (.A1(b[3]), .A2(a[3]), .ZN(n_45));
   OR2_X1 i_105 (.A1(b[4]), .A2(a[4]), .ZN(n_46));
   NAND3_X1 i_106 (.A1(n_50), .A2(n_49), .A3(n_48), .ZN(n_47));
   NAND2_X1 i_107 (.A1(b[2]), .A2(a[2]), .ZN(n_48));
   NAND2_X1 i_108 (.A1(b[3]), .A2(a[3]), .ZN(n_49));
   NAND3_X1 i_109 (.A1(n_53), .A2(n_51), .A3(n_52), .ZN(n_50));
   OR2_X1 i_110 (.A1(b[1]), .A2(a[1]), .ZN(n_51));
   OR2_X1 i_111 (.A1(b[2]), .A2(a[2]), .ZN(n_52));
   NAND2_X1 i_112 (.A1(n_15), .A2(n_22), .ZN(n_53));
   NAND2_X1 i_113 (.A1(b[9]), .A2(a[9]), .ZN(n_54));
   INV_X1 i_114 (.A(n_56), .ZN(n_55));
   NOR2_X1 i_115 (.A1(b[9]), .A2(a[9]), .ZN(n_56));
   INV_X1 i_116 (.A(a[8]), .ZN(n_57));
   INV_X1 i_117 (.A(b[8]), .ZN(n_58));
   AOI22_X1 i_118 (.A1(n_54), .A2(n_60), .B1(n_63), .B2(n_59), .ZN(p_0[10]));
   AND3_X1 i_119 (.A1(n_62), .A2(n_61), .A3(n_80), .ZN(n_59));
   AOI22_X1 i_120 (.A1(n_62), .A2(n_61), .B1(n_80), .B2(n_24), .ZN(n_60));
   OR2_X1 i_121 (.A1(a[10]), .A2(b[10]), .ZN(n_61));
   NAND2_X1 i_122 (.A1(a[10]), .A2(b[10]), .ZN(n_62));
   NAND3_X1 i_123 (.A1(n_29), .A2(n_54), .A3(n_25), .ZN(n_63));
   INV_X1 i_124 (.A(n_56), .ZN(n_80));
   NOR2_X1 i_125 (.A1(a[11]), .A2(b[11]), .ZN(n_81));
   INV_X1 i_126 (.A(n_81), .ZN(n_83));
   NAND2_X1 i_127 (.A1(a[11]), .A2(b[11]), .ZN(n_84));
   NAND3_X1 i_128 (.A1(n_61), .A2(n_80), .A3(n_63), .ZN(n_85));
   NAND2_X1 i_129 (.A1(n_85), .A2(n_62), .ZN(n_86));
   NAND2_X1 i_130 (.A1(n_83), .A2(n_84), .ZN(n_87));
   XNOR2_X1 i_131 (.A(n_86), .B(n_87), .ZN(p_0[11]));
   OAI21_X1 i_132 (.A(n_89), .B1(b[12]), .B2(a[12]), .ZN(n_88));
   NAND2_X1 i_133 (.A1(b[12]), .A2(a[12]), .ZN(n_89));
   NOR2_X1 i_134 (.A1(b[12]), .A2(a[12]), .ZN(n_90));
   NAND2_X1 i_135 (.A1(n_93), .A2(n_92), .ZN(n_91));
   NAND2_X1 i_136 (.A1(a[18]), .A2(b[18]), .ZN(n_92));
   OR2_X1 i_137 (.A1(a[18]), .A2(b[18]), .ZN(n_93));
   AOI21_X1 i_138 (.A(n_97), .B1(a[19]), .B2(b[19]), .ZN(n_94));
   NAND2_X1 i_139 (.A1(a[19]), .A2(b[19]), .ZN(n_95));
   INV_X1 i_140 (.A(n_97), .ZN(n_96));
   NOR2_X1 i_141 (.A1(a[19]), .A2(b[19]), .ZN(n_97));
   OAI21_X1 i_142 (.A(n_102), .B1(a[20]), .B2(b[20]), .ZN(n_101));
   NAND2_X1 i_143 (.A1(a[20]), .A2(b[20]), .ZN(n_102));
   NOR2_X1 i_144 (.A1(a[20]), .A2(b[20]), .ZN(n_103));
   NAND2_X1 i_145 (.A1(a[21]), .A2(b[21]), .ZN(n_104));
   NOR2_X1 i_146 (.A1(a[17]), .A2(b[17]), .ZN(n_105));
   INV_X1 i_147 (.A(n_105), .ZN(n_106));
   NAND2_X1 i_148 (.A1(a[16]), .A2(b[16]), .ZN(n_107));
   NAND2_X1 i_149 (.A1(a[17]), .A2(b[17]), .ZN(n_108));
   NAND2_X1 i_150 (.A1(a[15]), .A2(b[15]), .ZN(n_109));
   NAND2_X1 i_151 (.A1(a[14]), .A2(b[14]), .ZN(n_110));
   OR2_X1 i_152 (.A1(a[13]), .A2(b[13]), .ZN(n_111));
   NOR2_X1 i_153 (.A1(a[14]), .A2(b[14]), .ZN(n_112));
   INV_X1 i_154 (.A(n_112), .ZN(n_113));
   NOR2_X1 i_155 (.A1(a[15]), .A2(b[15]), .ZN(n_115));
   INV_X1 i_156 (.A(n_115), .ZN(n_116));
   NAND2_X1 i_157 (.A1(a[13]), .A2(b[13]), .ZN(n_117));
   INV_X1 i_158 (.A(n_31), .ZN(n_118));
   NAND3_X1 i_159 (.A1(n_55), .A2(n_83), .A3(n_61), .ZN(n_119));
   AOI211_X1 i_160 (.A(n_118), .B(n_119), .C1(n_57), .C2(n_58), .ZN(n_120));
   AOI21_X1 i_161 (.A(n_119), .B1(n_25), .B2(n_54), .ZN(n_121));
   INV_X1 i_162 (.A(n_84), .ZN(n_122));
   NOR2_X1 i_163 (.A1(n_81), .A2(n_62), .ZN(n_123));
   NOR4_X1 i_164 (.A1(n_120), .A2(n_121), .A3(n_122), .A4(n_123), .ZN(n_124));
   NAND3_X1 i_165 (.A1(n_116), .A2(n_111), .A3(n_113), .ZN(n_125));
   NOR3_X1 i_166 (.A1(n_124), .A2(n_90), .A3(n_125), .ZN(n_126));
   INV_X1 i_167 (.A(n_109), .ZN(n_127));
   NOR2_X1 i_168 (.A1(n_110), .A2(n_115), .ZN(n_128));
   AOI21_X1 i_169 (.A(n_125), .B1(n_89), .B2(n_117), .ZN(n_129));
   OR4_X1 i_170 (.A1(n_126), .A2(n_127), .A3(n_128), .A4(n_129), .ZN(n_130));
   INV_X1 i_171 (.A(a[16]), .ZN(n_131));
   INV_X1 i_172 (.A(b[16]), .ZN(n_132));
   NAND3_X1 i_173 (.A1(n_106), .A2(n_96), .A3(n_93), .ZN(n_133));
   AOI21_X1 i_174 (.A(n_133), .B1(n_107), .B2(n_108), .ZN(n_134));
   OAI21_X1 i_175 (.A(n_95), .B1(n_97), .B2(n_92), .ZN(n_135));
   AOI21_X1 i_176 (.A(n_133), .B1(n_131), .B2(n_132), .ZN(n_136));
   AOI211_X1 i_177 (.A(n_134), .B(n_135), .C1(n_130), .C2(n_136), .ZN(n_137));
   OAI211_X1 i_178 (.A(n_102), .B(n_104), .C1(n_137), .C2(n_103), .ZN(n_138));
   OR2_X1 i_179 (.A1(a[21]), .A2(b[21]), .ZN(n_139));
   NOR2_X1 i_180 (.A1(a[22]), .A2(b[22]), .ZN(n_140));
   NAND2_X1 i_181 (.A1(n_138), .A2(n_139), .ZN(n_141));
   INV_X1 i_182 (.A(n_140), .ZN(n_142));
   NAND2_X1 i_183 (.A1(a[22]), .A2(b[22]), .ZN(n_143));
   NAND2_X1 i_184 (.A1(n_142), .A2(n_143), .ZN(n_144));
   XOR2_X1 i_185 (.A(n_141), .B(n_144), .Z(p_0[22]));
   XNOR2_X1 i_186 (.A(n_146), .B(n_145), .ZN(p_0[23]));
   NAND2_X1 i_187 (.A1(n_149), .A2(n_148), .ZN(n_145));
   AOI21_X1 i_188 (.A(n_140), .B1(n_143), .B2(n_147), .ZN(n_146));
   NAND2_X1 i_189 (.A1(n_138), .A2(n_139), .ZN(n_147));
   NAND2_X1 i_190 (.A1(a[23]), .A2(b[23]), .ZN(n_148));
   INV_X1 i_191 (.A(n_150), .ZN(n_149));
   NOR2_X1 i_192 (.A1(a[23]), .A2(b[23]), .ZN(n_150));
   XNOR2_X1 i_193 (.A(n_152), .B(n_151), .ZN(p_0[24]));
   NAND2_X1 i_194 (.A1(n_161), .A2(n_160), .ZN(n_151));
   OAI21_X1 i_195 (.A(n_156), .B1(n_137), .B2(n_153), .ZN(n_152));
   INV_X1 i_196 (.A(n_154), .ZN(n_153));
   NOR2_X1 i_197 (.A1(n_103), .A2(n_159), .ZN(n_154));
   INV_X1 i_198 (.A(n_156), .ZN(n_155));
   NOR2_X1 i_199 (.A1(n_158), .A2(n_157), .ZN(n_156));
   OAI21_X1 i_200 (.A(n_148), .B1(n_150), .B2(n_143), .ZN(n_157));
   AOI21_X1 i_201 (.A(n_159), .B1(n_102), .B2(n_104), .ZN(n_158));
   NAND3_X1 i_202 (.A1(n_139), .A2(n_142), .A3(n_149), .ZN(n_159));
   NAND2_X1 i_203 (.A1(b[24]), .A2(a[24]), .ZN(n_160));
   NAND2_X1 i_204 (.A1(n_163), .A2(n_162), .ZN(n_161));
   INV_X1 i_205 (.A(a[24]), .ZN(n_162));
   INV_X1 i_206 (.A(b[24]), .ZN(n_163));
   OR2_X1 i_207 (.A1(a[25]), .A2(b[25]), .ZN(n_164));
   NAND2_X1 i_208 (.A1(n_152), .A2(n_161), .ZN(n_165));
   NAND2_X1 i_209 (.A1(a[25]), .A2(b[25]), .ZN(n_166));
   OR2_X1 i_210 (.A1(a[26]), .A2(b[26]), .ZN(n_167));
   NAND2_X1 i_211 (.A1(a[26]), .A2(b[26]), .ZN(n_168));
   NAND3_X1 i_212 (.A1(n_166), .A2(n_165), .A3(n_160), .ZN(n_169));
   NAND2_X1 i_213 (.A1(n_169), .A2(n_164), .ZN(n_170));
   NAND2_X1 i_214 (.A1(n_167), .A2(n_168), .ZN(n_171));
   XOR2_X1 i_215 (.A(n_170), .B(n_171), .Z(p_0[26]));
   XNOR2_X1 i_216 (.A(n_175), .B(n_172), .ZN(p_0[27]));
   OAI21_X1 i_218 (.A(n_168), .B1(n_174), .B2(n_173), .ZN(n_172));
   AND3_X1 i_219 (.A1(n_165), .A2(n_160), .A3(n_166), .ZN(n_173));
   NAND2_X1 i_220 (.A1(n_164), .A2(n_167), .ZN(n_174));
   NAND2_X1 i_221 (.A1(n_177), .A2(n_176), .ZN(n_175));
   NAND2_X1 i_222 (.A1(b[27]), .A2(a[27]), .ZN(n_176));
   INV_X1 i_223 (.A(n_178), .ZN(n_177));
   NOR2_X1 i_224 (.A1(b[27]), .A2(a[27]), .ZN(n_178));
   AND3_X1 i_225 (.A1(n_182), .A2(n_180), .A3(n_181), .ZN(n_179));
   NAND2_X1 i_226 (.A1(b[30]), .A2(a[30]), .ZN(n_180));
   NAND2_X1 i_227 (.A1(b[29]), .A2(a[29]), .ZN(n_181));
   INV_X1 i_228 (.A(n_183), .ZN(n_182));
   NOR2_X1 i_229 (.A1(b[29]), .A2(a[29]), .ZN(n_183));
   AOI211_X1 i_230 (.A(n_186), .B(n_185), .C1(n_155), .C2(n_187), .ZN(n_184));
   OAI21_X1 i_231 (.A(n_176), .B1(n_178), .B2(n_168), .ZN(n_185));
   AOI21_X1 i_232 (.A(n_188), .B1(n_160), .B2(n_166), .ZN(n_186));
   AOI21_X1 i_233 (.A(n_188), .B1(n_163), .B2(n_162), .ZN(n_187));
   NAND3_X1 i_234 (.A1(n_164), .A2(n_167), .A3(n_177), .ZN(n_188));
   NOR2_X1 i_235 (.A1(n_191), .A2(n_190), .ZN(n_189));
   OAI21_X1 i_236 (.A(n_211), .B1(n_180), .B2(n_209), .ZN(n_190));
   AOI21_X1 i_237 (.A(n_203), .B1(n_181), .B2(n_192), .ZN(n_191));
   NAND2_X1 i_238 (.A1(b[28]), .A2(a[28]), .ZN(n_192));
   NAND3_X1 i_239 (.A1(n_182), .A2(n_204), .A3(n_208), .ZN(n_203));
   INV_X1 i_240 (.A(n_207), .ZN(n_204));
   NOR2_X1 i_241 (.A1(b[30]), .A2(a[30]), .ZN(n_207));
   INV_X1 i_242 (.A(n_209), .ZN(n_208));
   NOR2_X1 i_243 (.A1(b[31]), .A2(a[31]), .ZN(n_209));
   NAND2_X1 i_244 (.A1(b[31]), .A2(a[31]), .ZN(n_211));
endmodule

module adderPlus(a, b, sum, cout);
   input [31:0]a;
   input [31:0]b;
   output [31:0]sum;
   output cout;

   datapath i_0 (.b(b), .a(a), .p_0({cout, sum[31], sum[30], sum[29], sum[28], 
      sum[27], sum[26], sum[25], sum[24], sum[23], sum[22], sum[21], sum[20], 
      sum[19], sum[18], sum[17], sum[16], sum[15], sum[14], sum[13], sum[12], 
      sum[11], sum[10], sum[9], sum[8], sum[7], sum[6], sum[5], sum[4], sum[3], 
      sum[2], sum[1], sum[0]}));
endmodule

module fullAdder__3_2(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   AND2_X1 i_0_1 (.A1(y), .A2(cin), .ZN(cout));
   XOR2_X1 i_0_0 (.A(cin), .B(y), .Z(sum));
endmodule

module fullAdder__3_5(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(y), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(x), .A2(cin), .ZN(n_0_2));
   OR2_X1 i_0_5 (.A1(x), .A2(cin), .ZN(n_0_3));
endmodule

module fullAdder__3_8(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_11(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_14(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_17(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_20(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_23(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_26(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_29(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_32(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_1;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
   XOR2_X1 i_0_2 (.A(y), .B(n_0_1), .Z(sum));
   XOR2_X1 i_0_3 (.A(cin), .B(x), .Z(n_0_1));
endmodule

module fullAdder__3_35(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_38(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_41(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_44(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_47(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_50(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_53(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_56(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_59(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_62(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_65(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_68(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_71(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_74(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_77(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_80(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_83(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_86(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__3_89(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module halfAdder(x, y, sum, cout);
   input x;
   input y;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(x), .A2(y), .ZN(cout));
endmodule

module PartialAdder(a, b, c, s1, c1);
   input [32:0]a;
   input [31:0]b;
   input [31:0]c;
   output [32:0]s1;
   output [31:0]c1;

   fullAdder__3_2 fa31 (.x(), .y(b[31]), .cin(c[30]), .sum(s1[31]), .cout(c1[31]));
   fullAdder__3_5 fa30 (.x(a[31]), .y(b[30]), .cin(c[29]), .sum(s1[30]), 
      .cout(c1[30]));
   fullAdder__3_8 fa29 (.x(a[30]), .y(b[29]), .cin(c[28]), .sum(s1[29]), 
      .cout(c1[29]));
   fullAdder__3_11 fa28 (.x(a[29]), .y(b[28]), .cin(c[27]), .sum(s1[28]), 
      .cout(c1[28]));
   fullAdder__3_14 fa27 (.x(a[28]), .y(b[27]), .cin(c[26]), .sum(s1[27]), 
      .cout(c1[27]));
   fullAdder__3_17 fa26 (.x(a[27]), .y(b[26]), .cin(c[25]), .sum(s1[26]), 
      .cout(c1[26]));
   fullAdder__3_20 fa25 (.x(a[26]), .y(b[25]), .cin(c[24]), .sum(s1[25]), 
      .cout(c1[25]));
   fullAdder__3_23 fa24 (.x(a[25]), .y(b[24]), .cin(c[23]), .sum(s1[24]), 
      .cout(c1[24]));
   fullAdder__3_26 fa23 (.x(a[24]), .y(b[23]), .cin(c[22]), .sum(s1[23]), 
      .cout(c1[23]));
   fullAdder__3_29 fa22 (.x(a[23]), .y(b[22]), .cin(c[21]), .sum(s1[22]), 
      .cout(c1[22]));
   fullAdder__3_32 fa21 (.x(a[22]), .y(b[21]), .cin(c[20]), .sum(s1[21]), 
      .cout(c1[21]));
   fullAdder__3_35 fa20 (.x(a[21]), .y(b[20]), .cin(c[19]), .sum(s1[20]), 
      .cout(c1[20]));
   fullAdder__3_38 fa19 (.x(a[20]), .y(b[19]), .cin(c[18]), .sum(s1[19]), 
      .cout(c1[19]));
   fullAdder__3_41 fa18 (.x(a[19]), .y(b[18]), .cin(c[17]), .sum(s1[18]), 
      .cout(c1[18]));
   fullAdder__3_44 fa17 (.x(a[18]), .y(b[17]), .cin(c[16]), .sum(s1[17]), 
      .cout(c1[17]));
   fullAdder__3_47 fa16 (.x(a[17]), .y(b[16]), .cin(c[15]), .sum(s1[16]), 
      .cout(c1[16]));
   fullAdder__3_50 fa15 (.x(a[16]), .y(b[15]), .cin(c[14]), .sum(s1[15]), 
      .cout(c1[15]));
   fullAdder__3_53 fa14 (.x(a[15]), .y(b[14]), .cin(c[13]), .sum(s1[14]), 
      .cout(c1[14]));
   fullAdder__3_56 fa13 (.x(a[14]), .y(b[13]), .cin(c[12]), .sum(s1[13]), 
      .cout(c1[13]));
   fullAdder__3_59 fa12 (.x(a[13]), .y(b[12]), .cin(c[11]), .sum(s1[12]), 
      .cout(c1[12]));
   fullAdder__3_62 fa11 (.x(a[12]), .y(b[11]), .cin(c[10]), .sum(s1[11]), 
      .cout(c1[11]));
   fullAdder__3_65 fa10 (.x(a[11]), .y(b[10]), .cin(c[9]), .sum(s1[10]), 
      .cout(c1[10]));
   fullAdder__3_68 fa9 (.x(a[10]), .y(b[9]), .cin(c[8]), .sum(s1[9]), .cout(
      c1[9]));
   fullAdder__3_71 fa8 (.x(a[9]), .y(b[8]), .cin(c[7]), .sum(s1[8]), .cout(c1[8]));
   fullAdder__3_74 fa7 (.x(a[8]), .y(b[7]), .cin(c[6]), .sum(s1[7]), .cout(c1[7]));
   fullAdder__3_77 fa6 (.x(a[7]), .y(b[6]), .cin(c[5]), .sum(s1[6]), .cout(c1[6]));
   fullAdder__3_80 fa5 (.x(a[6]), .y(b[5]), .cin(c[4]), .sum(s1[5]), .cout(c1[5]));
   fullAdder__3_83 fa4 (.x(a[5]), .y(b[4]), .cin(c[3]), .sum(s1[4]), .cout(c1[4]));
   fullAdder__3_86 fa3 (.x(a[4]), .y(b[3]), .cin(c[2]), .sum(s1[3]), .cout(c1[3]));
   fullAdder__3_89 fa2 (.x(a[3]), .y(b[2]), .cin(c[1]), .sum(s1[2]), .cout(c1[2]));
   fullAdder fa1 (.x(a[2]), .y(b[1]), .cin(c[0]), .sum(s1[1]), .cout(c1[1]));
   halfAdder ha1 (.x(a[1]), .y(b[0]), .sum(s1[0]), .cout(c1[0]));
endmodule

module datapath__0_4(p_0, b);
   output [31:0]p_0;
   input [31:0]b;

   XOR2_X1 i_0 (.A(b[1]), .B(b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(b[2]), .B1(b[1]), .B2(b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(b[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(b[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(b[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(b[6]), .B1(n_27), .B2(b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(b[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(b[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(b[9]), .B1(n_25), .B2(b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(b[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(b[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(b[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(b[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(b[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(b[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(b[16]), .B1(n_19), .B2(b[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(b[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(b[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(b[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(b[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(b[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(b[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(b[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(b[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(b[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(b[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(b[27]), .B1(n_9), .B2(b[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(b[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(b[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(b[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(b[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(b[28]), .A3(b[29]), .A4(b[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(b[28]), .A3(b[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(b[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(b[26]), .A3(b[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(b[23]), .A3(b[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(b[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(b[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(b[18]), .A3(b[19]), .A4(b[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(b[18]), .A3(b[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(b[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(b[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(b[15]), .A3(b[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(b[12]), .A3(b[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(b[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(b[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(b[8]), .A3(b[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(b[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(b[5]), .A3(b[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(b[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(b[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(b[2]), .A2(b[1]), .A3(b[0]), .ZN(n_29));
   INV_X1 i_61 (.A(b[11]), .ZN(n_30));
   INV_X1 i_62 (.A(b[14]), .ZN(n_31));
   INV_X1 i_63 (.A(b[21]), .ZN(n_32));
   INV_X1 i_64 (.A(b[25]), .ZN(n_33));
endmodule

module datapath__0_3(p_0, a);
   output [31:0]p_0;
   input [31:0]a;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[1]));
   NAND2_X1 i_1 (.A1(n_4), .A2(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(a[0]), .A2(a[1]), .ZN(n_1));
   INV_X1 i_3 (.A(n_2), .ZN(p_0[2]));
   NAND2_X1 i_4 (.A1(n_3), .A2(n_7), .ZN(n_2));
   NAND2_X1 i_5 (.A1(n_4), .A2(a[2]), .ZN(n_3));
   NAND2_X1 i_6 (.A1(n_142), .A2(n_143), .ZN(n_4));
   INV_X1 i_7 (.A(n_5), .ZN(p_0[3]));
   NAND2_X1 i_8 (.A1(n_6), .A2(n_141), .ZN(n_5));
   NAND2_X1 i_9 (.A1(n_7), .A2(a[3]), .ZN(n_6));
   NAND3_X1 i_10 (.A1(n_142), .A2(n_144), .A3(n_143), .ZN(n_7));
   INV_X1 i_11 (.A(n_8), .ZN(p_0[4]));
   NAND2_X1 i_12 (.A1(n_13), .A2(n_9), .ZN(n_8));
   NAND2_X1 i_13 (.A1(n_141), .A2(a[4]), .ZN(n_9));
   INV_X1 i_14 (.A(n_10), .ZN(p_0[5]));
   XNOR2_X1 i_15 (.A(n_15), .B(n_104), .ZN(n_10));
   INV_X1 i_16 (.A(n_11), .ZN(p_0[6]));
   NAND2_X1 i_17 (.A1(n_12), .A2(n_14), .ZN(n_11));
   OAI21_X1 i_18 (.A(a[6]), .B1(n_13), .B2(a[5]), .ZN(n_12));
   INV_X1 i_19 (.A(n_15), .ZN(n_13));
   XNOR2_X1 i_20 (.A(n_14), .B(n_125), .ZN(p_0[7]));
   NAND3_X1 i_21 (.A1(n_15), .A2(n_124), .A3(n_104), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_141), .A2(a[4]), .ZN(n_15));
   INV_X1 i_23 (.A(n_16), .ZN(p_0[8]));
   NAND2_X1 i_24 (.A1(n_20), .A2(n_17), .ZN(n_16));
   NAND2_X1 i_25 (.A1(n_40), .A2(a[8]), .ZN(n_17));
   INV_X1 i_26 (.A(n_18), .ZN(p_0[9]));
   NAND2_X1 i_27 (.A1(n_19), .A2(n_21), .ZN(n_18));
   NAND2_X1 i_28 (.A1(n_20), .A2(a[9]), .ZN(n_19));
   NAND2_X1 i_29 (.A1(n_39), .A2(n_128), .ZN(n_20));
   AOI21_X1 i_30 (.A(n_37), .B1(n_21), .B2(a[10]), .ZN(p_0[10]));
   NAND3_X1 i_31 (.A1(n_39), .A2(n_129), .A3(n_128), .ZN(n_21));
   INV_X1 i_32 (.A(n_22), .ZN(p_0[11]));
   NAND2_X1 i_33 (.A1(n_31), .A2(n_23), .ZN(n_22));
   NAND2_X1 i_34 (.A1(n_38), .A2(a[11]), .ZN(n_23));
   INV_X1 i_35 (.A(n_24), .ZN(p_0[12]));
   NAND2_X1 i_36 (.A1(n_25), .A2(n_28), .ZN(n_24));
   NAND2_X1 i_37 (.A1(n_31), .A2(a[12]), .ZN(n_25));
   INV_X1 i_38 (.A(n_26), .ZN(p_0[13]));
   OAI22_X1 i_39 (.A1(n_135), .A2(n_27), .B1(n_31), .B2(n_42), .ZN(n_26));
   INV_X1 i_40 (.A(n_28), .ZN(n_27));
   NAND3_X1 i_41 (.A1(n_37), .A2(n_134), .A3(n_133), .ZN(n_28));
   NOR2_X1 i_42 (.A1(n_29), .A2(n_35), .ZN(p_0[14]));
   AOI21_X1 i_43 (.A(n_138), .B1(n_30), .B2(n_41), .ZN(n_29));
   INV_X1 i_44 (.A(n_31), .ZN(n_30));
   NAND2_X1 i_45 (.A1(n_37), .A2(n_133), .ZN(n_31));
   INV_X1 i_46 (.A(n_32), .ZN(p_0[15]));
   OAI21_X1 i_47 (.A(n_33), .B1(n_35), .B2(n_139), .ZN(n_32));
   NAND4_X1 i_48 (.A1(n_37), .A2(n_133), .A3(n_34), .A4(n_41), .ZN(n_33));
   INV_X1 i_49 (.A(n_137), .ZN(n_34));
   INV_X1 i_50 (.A(n_36), .ZN(n_35));
   NAND4_X1 i_51 (.A1(n_37), .A2(n_138), .A3(n_133), .A4(n_41), .ZN(n_36));
   INV_X1 i_52 (.A(n_38), .ZN(n_37));
   NAND2_X1 i_53 (.A1(n_39), .A2(n_126), .ZN(n_38));
   INV_X1 i_54 (.A(n_40), .ZN(n_39));
   NAND2_X1 i_55 (.A1(n_140), .A2(n_120), .ZN(n_40));
   INV_X1 i_56 (.A(n_42), .ZN(n_41));
   NAND2_X1 i_57 (.A1(n_135), .A2(n_134), .ZN(n_42));
   INV_X1 i_58 (.A(n_43), .ZN(p_0[16]));
   XNOR2_X1 i_59 (.A(n_87), .B(a[16]), .ZN(n_43));
   INV_X1 i_60 (.A(n_44), .ZN(p_0[17]));
   NAND2_X1 i_61 (.A1(n_45), .A2(n_46), .ZN(n_44));
   OAI21_X1 i_62 (.A(a[17]), .B1(n_87), .B2(a[16]), .ZN(n_45));
   AOI21_X1 i_63 (.A(n_84), .B1(n_46), .B2(a[18]), .ZN(p_0[18]));
   NAND3_X1 i_64 (.A1(n_86), .A2(n_122), .A3(n_108), .ZN(n_46));
   INV_X1 i_65 (.A(n_47), .ZN(p_0[19]));
   NAND2_X1 i_66 (.A1(n_48), .A2(n_88), .ZN(n_47));
   NAND2_X1 i_67 (.A1(n_85), .A2(a[19]), .ZN(n_48));
   NOR2_X1 i_68 (.A1(n_49), .A2(n_51), .ZN(p_0[24]));
   NOR2_X1 i_69 (.A1(n_67), .A2(n_81), .ZN(n_49));
   INV_X1 i_70 (.A(n_50), .ZN(p_0[25]));
   OAI21_X1 i_71 (.A(n_55), .B1(n_51), .B2(n_82), .ZN(n_50));
   INV_X1 i_72 (.A(n_52), .ZN(n_51));
   NAND3_X1 i_73 (.A1(n_100), .A2(n_86), .A3(n_81), .ZN(n_52));
   INV_X1 i_74 (.A(n_53), .ZN(p_0[26]));
   NAND2_X1 i_75 (.A1(n_54), .A2(n_56), .ZN(n_53));
   NAND2_X1 i_76 (.A1(n_55), .A2(a[26]), .ZN(n_54));
   NAND3_X1 i_77 (.A1(n_100), .A2(n_86), .A3(n_57), .ZN(n_55));
   AOI21_X1 i_78 (.A(n_63), .B1(n_56), .B2(a[27]), .ZN(p_0[27]));
   NAND4_X1 i_79 (.A1(n_100), .A2(n_86), .A3(n_58), .A4(n_57), .ZN(n_56));
   INV_X1 i_80 (.A(n_80), .ZN(n_57));
   INV_X1 i_81 (.A(a[26]), .ZN(n_58));
   INV_X1 i_82 (.A(n_59), .ZN(p_0[28]));
   NAND2_X1 i_83 (.A1(n_60), .A2(n_61), .ZN(n_59));
   NAND2_X1 i_84 (.A1(n_64), .A2(a[28]), .ZN(n_60));
   AOI22_X1 i_85 (.A1(n_61), .A2(a[29]), .B1(n_63), .B2(n_73), .ZN(p_0[29]));
   NAND4_X1 i_86 (.A1(n_100), .A2(n_86), .A3(n_75), .A4(n_78), .ZN(n_61));
   AOI22_X1 i_87 (.A1(n_62), .A2(a[30]), .B1(n_63), .B2(n_71), .ZN(p_0[30]));
   NAND4_X1 i_88 (.A1(n_100), .A2(n_86), .A3(n_78), .A4(n_73), .ZN(n_62));
   INV_X1 i_89 (.A(n_64), .ZN(n_63));
   NAND3_X1 i_90 (.A1(n_100), .A2(n_86), .A3(n_78), .ZN(n_64));
   INV_X1 i_91 (.A(n_65), .ZN(p_0[31]));
   NAND2_X1 i_92 (.A1(n_66), .A2(n_69), .ZN(n_65));
   NAND4_X1 i_93 (.A1(n_67), .A2(n_68), .A3(n_78), .A4(n_71), .ZN(n_66));
   INV_X1 i_94 (.A(n_99), .ZN(n_67));
   INV_X1 i_95 (.A(a[31]), .ZN(n_68));
   NAND2_X1 i_96 (.A1(n_70), .A2(a[31]), .ZN(n_69));
   NAND4_X1 i_97 (.A1(n_100), .A2(n_86), .A3(n_78), .A4(n_71), .ZN(n_70));
   INV_X1 i_98 (.A(n_72), .ZN(n_71));
   NAND2_X1 i_99 (.A1(n_73), .A2(n_77), .ZN(n_72));
   INV_X1 i_100 (.A(n_74), .ZN(n_73));
   NAND2_X1 i_101 (.A1(n_76), .A2(n_75), .ZN(n_74));
   INV_X1 i_102 (.A(a[28]), .ZN(n_75));
   INV_X1 i_103 (.A(a[29]), .ZN(n_76));
   INV_X1 i_104 (.A(a[30]), .ZN(n_77));
   INV_X1 i_105 (.A(n_79), .ZN(n_78));
   OR3_X1 i_106 (.A1(n_80), .A2(a[27]), .A3(a[26]), .ZN(n_79));
   NAND2_X1 i_107 (.A1(n_82), .A2(n_81), .ZN(n_80));
   INV_X1 i_108 (.A(a[24]), .ZN(n_81));
   INV_X1 i_109 (.A(a[25]), .ZN(n_82));
   INV_X1 i_110 (.A(a[21]), .ZN(n_83));
   INV_X1 i_111 (.A(n_85), .ZN(n_84));
   NAND2_X1 i_112 (.A1(n_86), .A2(n_146), .ZN(n_85));
   INV_X1 i_113 (.A(n_87), .ZN(n_86));
   NAND2_X1 i_114 (.A1(n_118), .A2(n_140), .ZN(n_87));
   AOI21_X1 i_115 (.A(n_89), .B1(n_88), .B2(a[20]), .ZN(p_0[20]));
   NAND4_X1 i_116 (.A1(n_118), .A2(n_115), .A3(n_146), .A4(n_140), .ZN(n_88));
   INV_X1 i_117 (.A(n_90), .ZN(n_89));
   AOI21_X1 i_118 (.A(n_91), .B1(n_90), .B2(a[21]), .ZN(p_0[21]));
   NAND4_X1 i_119 (.A1(n_118), .A2(n_146), .A3(n_140), .A4(n_95), .ZN(n_90));
   INV_X1 i_120 (.A(n_92), .ZN(n_91));
   AOI21_X1 i_121 (.A(n_97), .B1(n_92), .B2(a[22]), .ZN(p_0[22]));
   NAND4_X1 i_122 (.A1(n_118), .A2(n_146), .A3(n_140), .A4(n_93), .ZN(n_92));
   INV_X1 i_123 (.A(n_94), .ZN(n_93));
   NAND2_X1 i_124 (.A1(n_95), .A2(n_83), .ZN(n_94));
   INV_X1 i_125 (.A(n_96), .ZN(n_95));
   NAND2_X1 i_126 (.A1(n_116), .A2(n_115), .ZN(n_96));
   INV_X1 i_127 (.A(n_112), .ZN(n_97));
   AOI21_X1 i_128 (.A(n_98), .B1(n_112), .B2(a[23]), .ZN(p_0[23]));
   INV_X1 i_129 (.A(n_99), .ZN(n_98));
   NAND4_X1 i_130 (.A1(n_100), .A2(n_105), .A3(n_140), .A4(n_111), .ZN(n_99));
   INV_X1 i_131 (.A(n_101), .ZN(n_100));
   NAND2_X1 i_132 (.A1(n_113), .A2(n_107), .ZN(n_101));
   INV_X1 i_133 (.A(n_106), .ZN(n_105));
   NAND3_X1 i_134 (.A1(n_126), .A2(n_109), .A3(n_102), .ZN(n_106));
   INV_X1 i_135 (.A(n_110), .ZN(n_109));
   NAND2_X1 i_136 (.A1(n_124), .A2(n_125), .ZN(n_110));
   NOR2_X1 i_142 (.A1(n_132), .A2(n_137), .ZN(n_111));
   NAND4_X1 i_143 (.A1(n_118), .A2(n_146), .A3(n_140), .A4(n_113), .ZN(n_112));
   INV_X1 i_137 (.A(n_114), .ZN(n_113));
   NAND4_X1 i_138 (.A1(n_83), .A2(n_116), .A3(n_115), .A4(n_117), .ZN(n_114));
   INV_X1 i_139 (.A(a[19]), .ZN(n_115));
   INV_X1 i_140 (.A(a[20]), .ZN(n_116));
   INV_X1 i_141 (.A(a[22]), .ZN(n_117));
   INV_X1 i_144 (.A(n_119), .ZN(n_118));
   NAND4_X1 i_145 (.A1(n_120), .A2(n_136), .A3(n_131), .A4(n_126), .ZN(n_119));
   INV_X1 i_146 (.A(n_121), .ZN(n_120));
   NAND4_X1 i_147 (.A1(n_103), .A2(n_104), .A3(n_124), .A4(n_125), .ZN(n_121));
   INV_X1 i_148 (.A(a[6]), .ZN(n_124));
   INV_X1 i_149 (.A(a[7]), .ZN(n_125));
   INV_X1 i_150 (.A(n_127), .ZN(n_126));
   NAND3_X1 i_151 (.A1(n_130), .A2(n_129), .A3(n_128), .ZN(n_127));
   INV_X1 i_152 (.A(a[8]), .ZN(n_128));
   INV_X1 i_153 (.A(a[9]), .ZN(n_129));
   INV_X1 i_154 (.A(a[10]), .ZN(n_130));
   INV_X1 i_155 (.A(n_132), .ZN(n_131));
   NAND3_X1 i_156 (.A1(n_134), .A2(n_133), .A3(n_135), .ZN(n_132));
   INV_X1 i_157 (.A(a[11]), .ZN(n_133));
   INV_X1 i_158 (.A(a[12]), .ZN(n_134));
   INV_X1 i_159 (.A(a[13]), .ZN(n_135));
   INV_X1 i_160 (.A(n_137), .ZN(n_136));
   NAND2_X1 i_161 (.A1(n_139), .A2(n_138), .ZN(n_137));
   INV_X1 i_162 (.A(a[14]), .ZN(n_138));
   INV_X1 i_163 (.A(a[15]), .ZN(n_139));
   INV_X1 i_164 (.A(n_141), .ZN(n_140));
   NAND4_X1 i_165 (.A1(n_142), .A2(n_145), .A3(n_144), .A4(n_143), .ZN(n_141));
   INV_X1 i_173 (.A(a[0]), .ZN(n_142));
   INV_X1 i_166 (.A(a[1]), .ZN(n_143));
   INV_X1 i_167 (.A(a[2]), .ZN(n_144));
   INV_X1 i_168 (.A(a[3]), .ZN(n_145));
   INV_X1 i_177 (.A(n_147), .ZN(n_146));
   NAND3_X1 i_178 (.A1(n_108), .A2(n_123), .A3(n_122), .ZN(n_147));
   NOR2_X1 i_169 (.A1(a[5]), .A2(a[4]), .ZN(n_102));
   INV_X1 i_170 (.A(a[4]), .ZN(n_103));
   INV_X1 i_171 (.A(a[5]), .ZN(n_104));
   NOR4_X1 i_172 (.A1(a[18]), .A2(a[16]), .A3(a[17]), .A4(a[23]), .ZN(n_107));
   INV_X1 i_174 (.A(a[16]), .ZN(n_108));
   INV_X1 i_175 (.A(a[17]), .ZN(n_122));
   INV_X1 i_176 (.A(a[18]), .ZN(n_123));
endmodule

module datapath__0_38(p_0, sum1);
   output [63:0]p_0;
   input [63:0]sum1;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[1]));
   XNOR2_X1 i_1 (.A(sum1[1]), .B(sum1[0]), .ZN(n_0));
   INV_X1 i_2 (.A(n_1), .ZN(p_0[2]));
   NAND2_X1 i_3 (.A1(n_173), .A2(n_2), .ZN(n_1));
   NAND2_X1 i_4 (.A1(sum1[2]), .A2(n_175), .ZN(n_2));
   INV_X1 i_5 (.A(n_3), .ZN(p_0[3]));
   NAND2_X1 i_6 (.A1(n_171), .A2(n_4), .ZN(n_3));
   NAND2_X1 i_7 (.A1(sum1[3]), .A2(n_173), .ZN(n_4));
   INV_X1 i_8 (.A(n_5), .ZN(p_0[4]));
   NAND2_X1 i_9 (.A1(n_169), .A2(n_6), .ZN(n_5));
   NAND2_X1 i_10 (.A1(sum1[4]), .A2(n_171), .ZN(n_6));
   INV_X1 i_11 (.A(n_7), .ZN(p_0[5]));
   NAND2_X1 i_12 (.A1(n_167), .A2(n_8), .ZN(n_7));
   NAND2_X1 i_13 (.A1(sum1[5]), .A2(n_169), .ZN(n_8));
   INV_X1 i_14 (.A(n_9), .ZN(p_0[6]));
   NAND2_X1 i_15 (.A1(n_165), .A2(n_10), .ZN(n_9));
   NAND2_X1 i_16 (.A1(sum1[6]), .A2(n_167), .ZN(n_10));
   INV_X1 i_17 (.A(n_11), .ZN(p_0[7]));
   NAND2_X1 i_18 (.A1(n_163), .A2(n_12), .ZN(n_11));
   NAND2_X1 i_19 (.A1(sum1[7]), .A2(n_165), .ZN(n_12));
   INV_X1 i_20 (.A(n_13), .ZN(p_0[8]));
   NAND2_X1 i_21 (.A1(n_161), .A2(n_14), .ZN(n_13));
   NAND2_X1 i_22 (.A1(sum1[8]), .A2(n_163), .ZN(n_14));
   INV_X1 i_23 (.A(n_15), .ZN(p_0[9]));
   NAND2_X1 i_24 (.A1(n_159), .A2(n_16), .ZN(n_15));
   NAND2_X1 i_25 (.A1(sum1[9]), .A2(n_161), .ZN(n_16));
   INV_X1 i_26 (.A(n_17), .ZN(p_0[10]));
   NAND2_X1 i_27 (.A1(n_157), .A2(n_18), .ZN(n_17));
   NAND2_X1 i_28 (.A1(sum1[10]), .A2(n_159), .ZN(n_18));
   INV_X1 i_29 (.A(n_19), .ZN(p_0[11]));
   NAND2_X1 i_30 (.A1(n_155), .A2(n_20), .ZN(n_19));
   NAND2_X1 i_31 (.A1(sum1[11]), .A2(n_157), .ZN(n_20));
   INV_X1 i_32 (.A(n_21), .ZN(p_0[12]));
   NAND2_X1 i_33 (.A1(n_153), .A2(n_22), .ZN(n_21));
   NAND2_X1 i_34 (.A1(sum1[12]), .A2(n_155), .ZN(n_22));
   INV_X1 i_35 (.A(n_23), .ZN(p_0[13]));
   NAND2_X1 i_36 (.A1(n_151), .A2(n_24), .ZN(n_23));
   NAND2_X1 i_37 (.A1(sum1[13]), .A2(n_153), .ZN(n_24));
   INV_X1 i_38 (.A(n_25), .ZN(p_0[14]));
   NAND2_X1 i_39 (.A1(n_149), .A2(n_26), .ZN(n_25));
   NAND2_X1 i_40 (.A1(sum1[14]), .A2(n_151), .ZN(n_26));
   INV_X1 i_41 (.A(n_27), .ZN(p_0[15]));
   NAND2_X1 i_42 (.A1(n_147), .A2(n_28), .ZN(n_27));
   NAND2_X1 i_43 (.A1(sum1[15]), .A2(n_149), .ZN(n_28));
   INV_X1 i_44 (.A(n_29), .ZN(p_0[16]));
   NAND2_X1 i_45 (.A1(n_145), .A2(n_30), .ZN(n_29));
   NAND2_X1 i_46 (.A1(sum1[16]), .A2(n_147), .ZN(n_30));
   INV_X1 i_47 (.A(n_31), .ZN(p_0[17]));
   NAND2_X1 i_48 (.A1(n_143), .A2(n_32), .ZN(n_31));
   NAND2_X1 i_49 (.A1(sum1[17]), .A2(n_145), .ZN(n_32));
   INV_X1 i_50 (.A(n_33), .ZN(p_0[18]));
   NAND2_X1 i_51 (.A1(n_141), .A2(n_34), .ZN(n_33));
   NAND2_X1 i_52 (.A1(sum1[18]), .A2(n_143), .ZN(n_34));
   INV_X1 i_53 (.A(n_35), .ZN(p_0[19]));
   NAND2_X1 i_54 (.A1(n_139), .A2(n_36), .ZN(n_35));
   NAND2_X1 i_55 (.A1(sum1[19]), .A2(n_141), .ZN(n_36));
   INV_X1 i_56 (.A(n_37), .ZN(p_0[20]));
   NAND2_X1 i_57 (.A1(n_137), .A2(n_38), .ZN(n_37));
   NAND2_X1 i_58 (.A1(sum1[20]), .A2(n_139), .ZN(n_38));
   INV_X1 i_59 (.A(n_39), .ZN(p_0[21]));
   NAND2_X1 i_60 (.A1(n_135), .A2(n_40), .ZN(n_39));
   NAND2_X1 i_61 (.A1(sum1[21]), .A2(n_137), .ZN(n_40));
   INV_X1 i_62 (.A(n_41), .ZN(p_0[22]));
   NAND2_X1 i_63 (.A1(n_224), .A2(n_42), .ZN(n_41));
   NAND2_X1 i_64 (.A1(sum1[22]), .A2(n_135), .ZN(n_42));
   INV_X1 i_65 (.A(n_43), .ZN(p_0[23]));
   NAND2_X1 i_66 (.A1(n_223), .A2(n_44), .ZN(n_43));
   NAND2_X1 i_67 (.A1(sum1[23]), .A2(n_224), .ZN(n_44));
   INV_X1 i_68 (.A(n_45), .ZN(p_0[24]));
   NAND2_X1 i_69 (.A1(n_221), .A2(n_46), .ZN(n_45));
   NAND2_X1 i_70 (.A1(sum1[24]), .A2(n_223), .ZN(n_46));
   INV_X1 i_71 (.A(n_47), .ZN(p_0[25]));
   NAND2_X1 i_72 (.A1(n_219), .A2(n_48), .ZN(n_47));
   NAND2_X1 i_73 (.A1(sum1[25]), .A2(n_221), .ZN(n_48));
   INV_X1 i_74 (.A(n_49), .ZN(p_0[26]));
   NAND2_X1 i_75 (.A1(n_218), .A2(n_50), .ZN(n_49));
   NAND2_X1 i_76 (.A1(sum1[26]), .A2(n_219), .ZN(n_50));
   INV_X1 i_77 (.A(n_51), .ZN(p_0[27]));
   NAND2_X1 i_78 (.A1(n_216), .A2(n_52), .ZN(n_51));
   NAND2_X1 i_79 (.A1(sum1[27]), .A2(n_218), .ZN(n_52));
   INV_X1 i_80 (.A(n_53), .ZN(p_0[28]));
   NAND2_X1 i_81 (.A1(n_215), .A2(n_54), .ZN(n_53));
   NAND2_X1 i_82 (.A1(n_216), .A2(sum1[28]), .ZN(n_54));
   INV_X1 i_83 (.A(n_55), .ZN(p_0[29]));
   NAND2_X1 i_84 (.A1(n_214), .A2(n_56), .ZN(n_55));
   NAND2_X1 i_85 (.A1(sum1[29]), .A2(n_215), .ZN(n_56));
   INV_X1 i_86 (.A(n_57), .ZN(p_0[30]));
   XNOR2_X1 i_87 (.A(sum1[30]), .B(n_214), .ZN(n_57));
   INV_X1 i_88 (.A(n_58), .ZN(p_0[31]));
   XNOR2_X1 i_89 (.A(n_213), .B(n_225), .ZN(n_58));
   INV_X1 i_90 (.A(n_59), .ZN(p_0[32]));
   XNOR2_X1 i_91 (.A(sum1[32]), .B(n_212), .ZN(n_59));
   INV_X1 i_92 (.A(n_60), .ZN(p_0[33]));
   XNOR2_X1 i_93 (.A(n_211), .B(n_226), .ZN(n_60));
   INV_X1 i_94 (.A(n_61), .ZN(p_0[34]));
   NAND2_X1 i_95 (.A1(n_209), .A2(n_62), .ZN(n_61));
   NAND2_X1 i_96 (.A1(n_210), .A2(sum1[34]), .ZN(n_62));
   INV_X1 i_97 (.A(n_63), .ZN(p_0[35]));
   NAND2_X1 i_98 (.A1(n_190), .A2(n_64), .ZN(n_63));
   NAND2_X1 i_99 (.A1(n_209), .A2(sum1[35]), .ZN(n_64));
   INV_X1 i_100 (.A(n_65), .ZN(p_0[36]));
   NAND2_X1 i_101 (.A1(n_208), .A2(n_66), .ZN(n_65));
   NAND2_X1 i_102 (.A1(n_190), .A2(sum1[36]), .ZN(n_66));
   INV_X1 i_103 (.A(n_67), .ZN(p_0[37]));
   NAND2_X1 i_104 (.A1(n_71), .A2(n_68), .ZN(n_67));
   NAND2_X1 i_105 (.A1(n_208), .A2(sum1[37]), .ZN(n_68));
   INV_X1 i_106 (.A(n_69), .ZN(p_0[38]));
   OAI21_X1 i_107 (.A(n_74), .B1(n_189), .B2(n_70), .ZN(n_69));
   INV_X1 i_108 (.A(n_71), .ZN(n_70));
   NAND2_X1 i_109 (.A1(n_207), .A2(n_228), .ZN(n_71));
   INV_X1 i_110 (.A(n_72), .ZN(p_0[39]));
   NAND2_X1 i_111 (.A1(n_73), .A2(n_206), .ZN(n_72));
   NAND2_X1 i_112 (.A1(n_74), .A2(sum1[39]), .ZN(n_73));
   NAND3_X1 i_113 (.A1(n_207), .A2(n_189), .A3(n_228), .ZN(n_74));
   INV_X1 i_114 (.A(n_75), .ZN(p_0[40]));
   XNOR2_X1 i_115 (.A(sum1[40]), .B(n_206), .ZN(n_75));
   INV_X1 i_116 (.A(n_76), .ZN(p_0[41]));
   XNOR2_X1 i_117 (.A(n_205), .B(n_229), .ZN(n_76));
   INV_X1 i_118 (.A(n_77), .ZN(p_0[42]));
   XNOR2_X1 i_119 (.A(n_204), .B(sum1[42]), .ZN(n_77));
   INV_X1 i_120 (.A(n_78), .ZN(p_0[43]));
   XNOR2_X1 i_121 (.A(n_187), .B(n_231), .ZN(n_78));
   INV_X1 i_122 (.A(n_79), .ZN(p_0[44]));
   NAND2_X1 i_123 (.A1(n_85), .A2(n_80), .ZN(n_79));
   NAND2_X1 i_124 (.A1(n_202), .A2(sum1[44]), .ZN(n_80));
   INV_X1 i_125 (.A(n_81), .ZN(p_0[45]));
   XNOR2_X1 i_126 (.A(n_185), .B(n_184), .ZN(n_81));
   INV_X1 i_127 (.A(n_82), .ZN(p_0[46]));
   XNOR2_X1 i_128 (.A(n_84), .B(n_233), .ZN(n_82));
   NOR2_X1 i_129 (.A1(n_83), .A2(n_199), .ZN(p_0[47]));
   AOI21_X1 i_130 (.A(n_183), .B1(n_84), .B2(n_233), .ZN(n_83));
   NOR2_X1 i_131 (.A1(n_85), .A2(sum1[45]), .ZN(n_84));
   INV_X1 i_132 (.A(n_185), .ZN(n_85));
   INV_X1 i_133 (.A(n_86), .ZN(p_0[48]));
   NAND2_X1 i_134 (.A1(n_92), .A2(n_87), .ZN(n_86));
   NAND2_X1 i_135 (.A1(n_200), .A2(sum1[48]), .ZN(n_87));
   INV_X1 i_136 (.A(n_88), .ZN(p_0[49]));
   XNOR2_X1 i_137 (.A(n_92), .B(sum1[49]), .ZN(n_88));
   AND2_X1 i_138 (.A1(n_89), .A2(n_90), .ZN(p_0[50]));
   OAI21_X1 i_139 (.A(sum1[50]), .B1(n_92), .B2(sum1[49]), .ZN(n_89));
   XNOR2_X1 i_140 (.A(n_90), .B(n_133), .ZN(p_0[51]));
   NAND3_X1 i_141 (.A1(n_91), .A2(n_132), .A3(n_131), .ZN(n_90));
   INV_X1 i_142 (.A(n_92), .ZN(n_91));
   NAND2_X1 i_143 (.A1(n_199), .A2(n_130), .ZN(n_92));
   INV_X1 i_144 (.A(n_93), .ZN(p_0[52]));
   NAND2_X1 i_145 (.A1(n_97), .A2(n_94), .ZN(n_93));
   NAND2_X1 i_146 (.A1(n_102), .A2(sum1[52]), .ZN(n_94));
   INV_X1 i_147 (.A(n_95), .ZN(p_0[53]));
   NAND2_X1 i_148 (.A1(n_96), .A2(n_100), .ZN(n_95));
   NAND2_X1 i_149 (.A1(n_97), .A2(sum1[53]), .ZN(n_96));
   NAND2_X1 i_150 (.A1(n_101), .A2(n_127), .ZN(n_97));
   INV_X1 i_151 (.A(n_98), .ZN(p_0[54]));
   XNOR2_X1 i_152 (.A(n_100), .B(sum1[54]), .ZN(n_98));
   AOI21_X1 i_153 (.A(n_181), .B1(n_99), .B2(sum1[55]), .ZN(p_0[55]));
   OR2_X1 i_154 (.A1(n_100), .A2(sum1[54]), .ZN(n_99));
   NAND3_X1 i_155 (.A1(n_101), .A2(n_128), .A3(n_127), .ZN(n_100));
   INV_X1 i_156 (.A(n_102), .ZN(n_101));
   NAND2_X1 i_157 (.A1(n_199), .A2(n_234), .ZN(n_102));
   INV_X1 i_158 (.A(n_103), .ZN(p_0[56]));
   NAND2_X1 i_159 (.A1(n_107), .A2(n_104), .ZN(n_103));
   NAND2_X1 i_160 (.A1(n_182), .A2(sum1[56]), .ZN(n_104));
   INV_X1 i_161 (.A(n_105), .ZN(p_0[57]));
   OAI21_X1 i_162 (.A(n_110), .B1(n_106), .B2(n_237), .ZN(n_105));
   INV_X1 i_163 (.A(n_107), .ZN(n_106));
   NAND2_X1 i_164 (.A1(n_181), .A2(n_236), .ZN(n_107));
   INV_X1 i_165 (.A(n_108), .ZN(p_0[58]));
   NAND2_X1 i_166 (.A1(n_109), .A2(n_180), .ZN(n_108));
   NAND2_X1 i_167 (.A1(n_110), .A2(sum1[58]), .ZN(n_109));
   NAND2_X1 i_168 (.A1(n_124), .A2(n_181), .ZN(n_110));
   INV_X1 i_169 (.A(n_111), .ZN(p_0[59]));
   NAND2_X1 i_170 (.A1(n_123), .A2(n_112), .ZN(n_111));
   NAND2_X1 i_171 (.A1(n_180), .A2(sum1[59]), .ZN(n_112));
   NOR2_X1 i_172 (.A1(n_113), .A2(n_118), .ZN(p_0[60]));
   NOR2_X1 i_173 (.A1(n_122), .A2(n_179), .ZN(n_113));
   INV_X1 i_174 (.A(n_114), .ZN(p_0[62]));
   NAND2_X1 i_175 (.A1(n_115), .A2(n_121), .ZN(n_114));
   OAI21_X1 i_176 (.A(sum1[62]), .B1(n_195), .B2(sum1[61]), .ZN(n_115));
   INV_X1 i_177 (.A(n_116), .ZN(p_0[63]));
   NAND2_X1 i_178 (.A1(n_120), .A2(n_117), .ZN(n_116));
   NAND4_X1 i_179 (.A1(n_118), .A2(n_119), .A3(n_177), .A4(n_176), .ZN(n_117));
   INV_X1 i_180 (.A(n_195), .ZN(n_118));
   INV_X1 i_181 (.A(sum1[63]), .ZN(n_119));
   NAND2_X1 i_182 (.A1(n_121), .A2(sum1[63]), .ZN(n_120));
   NAND4_X1 i_183 (.A1(n_122), .A2(n_177), .A3(n_176), .A4(n_179), .ZN(n_121));
   INV_X1 i_184 (.A(n_123), .ZN(n_122));
   NAND4_X1 i_185 (.A1(n_124), .A2(n_178), .A3(n_238), .A4(n_181), .ZN(n_123));
   NOR2_X1 i_186 (.A1(sum1[57]), .A2(sum1[56]), .ZN(n_124));
   NAND3_X1 i_187 (.A1(n_128), .A2(n_127), .A3(n_126), .ZN(n_125));
   NOR2_X1 i_188 (.A1(sum1[54]), .A2(sum1[55]), .ZN(n_126));
   INV_X1 i_189 (.A(sum1[52]), .ZN(n_127));
   INV_X1 i_190 (.A(sum1[53]), .ZN(n_128));
   NAND4_X1 i_191 (.A1(n_132), .A2(n_131), .A3(n_133), .A4(n_130), .ZN(n_129));
   INV_X1 i_192 (.A(sum1[48]), .ZN(n_130));
   INV_X1 i_193 (.A(sum1[49]), .ZN(n_131));
   INV_X1 i_194 (.A(sum1[50]), .ZN(n_132));
   INV_X1 i_195 (.A(sum1[51]), .ZN(n_133));
   NOR2_X1 i_196 (.A1(sum1[22]), .A2(n_135), .ZN(n_134));
   INV_X1 i_197 (.A(n_136), .ZN(n_135));
   NOR2_X1 i_198 (.A1(sum1[21]), .A2(n_137), .ZN(n_136));
   INV_X1 i_199 (.A(n_138), .ZN(n_137));
   NOR2_X1 i_200 (.A1(sum1[20]), .A2(n_139), .ZN(n_138));
   INV_X1 i_201 (.A(n_140), .ZN(n_139));
   NOR2_X1 i_202 (.A1(sum1[19]), .A2(n_141), .ZN(n_140));
   INV_X1 i_203 (.A(n_142), .ZN(n_141));
   NOR2_X1 i_204 (.A1(sum1[18]), .A2(n_143), .ZN(n_142));
   INV_X1 i_205 (.A(n_144), .ZN(n_143));
   NOR2_X1 i_206 (.A1(sum1[17]), .A2(n_145), .ZN(n_144));
   INV_X1 i_207 (.A(n_146), .ZN(n_145));
   NOR2_X1 i_208 (.A1(sum1[16]), .A2(n_147), .ZN(n_146));
   INV_X1 i_209 (.A(n_148), .ZN(n_147));
   NOR2_X1 i_210 (.A1(sum1[15]), .A2(n_149), .ZN(n_148));
   INV_X1 i_211 (.A(n_150), .ZN(n_149));
   NOR2_X1 i_212 (.A1(sum1[14]), .A2(n_151), .ZN(n_150));
   INV_X1 i_213 (.A(n_152), .ZN(n_151));
   NOR2_X1 i_214 (.A1(sum1[13]), .A2(n_153), .ZN(n_152));
   INV_X1 i_215 (.A(n_154), .ZN(n_153));
   NOR2_X1 i_216 (.A1(sum1[12]), .A2(n_155), .ZN(n_154));
   INV_X1 i_217 (.A(n_156), .ZN(n_155));
   NOR2_X1 i_218 (.A1(sum1[11]), .A2(n_157), .ZN(n_156));
   INV_X1 i_219 (.A(n_158), .ZN(n_157));
   NOR2_X1 i_220 (.A1(sum1[10]), .A2(n_159), .ZN(n_158));
   INV_X1 i_221 (.A(n_160), .ZN(n_159));
   NOR2_X1 i_222 (.A1(sum1[9]), .A2(n_161), .ZN(n_160));
   INV_X1 i_223 (.A(n_162), .ZN(n_161));
   NOR2_X1 i_224 (.A1(sum1[8]), .A2(n_163), .ZN(n_162));
   INV_X1 i_225 (.A(n_164), .ZN(n_163));
   NOR2_X1 i_226 (.A1(sum1[7]), .A2(n_165), .ZN(n_164));
   INV_X1 i_227 (.A(n_166), .ZN(n_165));
   NOR2_X1 i_228 (.A1(sum1[6]), .A2(n_167), .ZN(n_166));
   INV_X1 i_229 (.A(n_168), .ZN(n_167));
   NOR2_X1 i_230 (.A1(sum1[5]), .A2(n_169), .ZN(n_168));
   INV_X1 i_231 (.A(n_170), .ZN(n_169));
   NOR2_X1 i_232 (.A1(sum1[4]), .A2(n_171), .ZN(n_170));
   INV_X1 i_233 (.A(n_172), .ZN(n_171));
   NOR2_X1 i_234 (.A1(sum1[3]), .A2(n_173), .ZN(n_172));
   INV_X1 i_235 (.A(n_174), .ZN(n_173));
   NOR2_X1 i_236 (.A1(sum1[2]), .A2(n_175), .ZN(n_174));
   OR2_X1 i_237 (.A1(sum1[1]), .A2(sum1[0]), .ZN(n_175));
   INV_X1 i_238 (.A(sum1[61]), .ZN(n_176));
   INV_X1 i_239 (.A(sum1[62]), .ZN(n_177));
   INV_X1 i_240 (.A(sum1[59]), .ZN(n_178));
   INV_X1 i_241 (.A(sum1[60]), .ZN(n_179));
   NAND3_X1 i_242 (.A1(n_197), .A2(n_238), .A3(n_237), .ZN(n_180));
   INV_X1 i_243 (.A(n_182), .ZN(n_181));
   NAND3_X1 i_244 (.A1(n_235), .A2(n_234), .A3(n_199), .ZN(n_182));
   INV_X1 i_245 (.A(sum1[47]), .ZN(n_183));
   INV_X1 i_246 (.A(sum1[45]), .ZN(n_184));
   INV_X1 i_247 (.A(n_186), .ZN(n_185));
   OR2_X1 i_248 (.A1(n_202), .A2(sum1[44]), .ZN(n_186));
   INV_X1 i_249 (.A(n_188), .ZN(n_187));
   NAND2_X1 i_250 (.A1(n_203), .A2(n_230), .ZN(n_188));
   INV_X1 i_251 (.A(sum1[38]), .ZN(n_189));
   OR2_X1 i_252 (.A1(n_209), .A2(sum1[35]), .ZN(n_190));
   INV_X1 i_253 (.A(n_191), .ZN(p_0[61]));
   NAND2_X1 i_254 (.A1(n_193), .A2(n_192), .ZN(n_191));
   NAND2_X1 i_255 (.A1(sum1[61]), .A2(n_195), .ZN(n_192));
   NAND2_X1 i_256 (.A1(n_239), .A2(n_194), .ZN(n_193));
   INV_X1 i_257 (.A(n_195), .ZN(n_194));
   NAND4_X1 i_258 (.A1(n_196), .A2(n_197), .A3(n_238), .A4(n_237), .ZN(n_195));
   NOR2_X1 i_259 (.A1(sum1[59]), .A2(sum1[60]), .ZN(n_196));
   INV_X1 i_260 (.A(n_198), .ZN(n_197));
   NAND4_X1 i_261 (.A1(n_235), .A2(n_234), .A3(n_236), .A4(n_199), .ZN(n_198));
   INV_X1 i_262 (.A(n_200), .ZN(n_199));
   NAND3_X1 i_263 (.A1(n_233), .A2(n_232), .A3(n_201), .ZN(n_200));
   INV_X1 i_264 (.A(n_202), .ZN(n_201));
   NAND3_X1 i_265 (.A1(n_203), .A2(n_231), .A3(n_230), .ZN(n_202));
   INV_X1 i_266 (.A(n_204), .ZN(n_203));
   NAND2_X1 i_267 (.A1(n_205), .A2(n_229), .ZN(n_204));
   NOR2_X1 i_268 (.A1(n_206), .A2(sum1[40]), .ZN(n_205));
   NAND3_X1 i_269 (.A1(n_207), .A2(n_228), .A3(n_227), .ZN(n_206));
   INV_X1 i_270 (.A(n_208), .ZN(n_207));
   OR3_X1 i_271 (.A1(n_209), .A2(sum1[35]), .A3(sum1[36]), .ZN(n_208));
   OR2_X1 i_272 (.A1(sum1[34]), .A2(n_210), .ZN(n_209));
   NAND2_X1 i_273 (.A1(n_211), .A2(n_226), .ZN(n_210));
   NOR2_X1 i_274 (.A1(sum1[32]), .A2(n_212), .ZN(n_211));
   NAND2_X1 i_275 (.A1(n_225), .A2(n_213), .ZN(n_212));
   NOR2_X1 i_276 (.A1(n_214), .A2(sum1[30]), .ZN(n_213));
   OR2_X1 i_277 (.A1(n_215), .A2(sum1[29]), .ZN(n_214));
   OR2_X1 i_278 (.A1(n_216), .A2(sum1[28]), .ZN(n_215));
   INV_X1 i_279 (.A(n_217), .ZN(n_216));
   NOR2_X1 i_280 (.A1(sum1[27]), .A2(n_218), .ZN(n_217));
   OR2_X1 i_281 (.A1(sum1[26]), .A2(n_219), .ZN(n_218));
   INV_X1 i_282 (.A(n_220), .ZN(n_219));
   NOR2_X1 i_283 (.A1(sum1[25]), .A2(n_221), .ZN(n_220));
   INV_X1 i_284 (.A(n_222), .ZN(n_221));
   NOR2_X1 i_285 (.A1(n_223), .A2(sum1[24]), .ZN(n_222));
   OR2_X1 i_286 (.A1(sum1[23]), .A2(n_224), .ZN(n_223));
   INV_X1 i_287 (.A(n_134), .ZN(n_224));
   INV_X1 i_288 (.A(sum1[31]), .ZN(n_225));
   INV_X1 i_289 (.A(sum1[33]), .ZN(n_226));
   NOR2_X1 i_290 (.A1(sum1[39]), .A2(sum1[38]), .ZN(n_227));
   INV_X1 i_291 (.A(sum1[37]), .ZN(n_228));
   INV_X1 i_292 (.A(sum1[41]), .ZN(n_229));
   INV_X1 i_293 (.A(sum1[42]), .ZN(n_230));
   INV_X1 i_294 (.A(sum1[43]), .ZN(n_231));
   NOR3_X1 i_295 (.A1(sum1[45]), .A2(sum1[47]), .A3(sum1[44]), .ZN(n_232));
   INV_X1 i_296 (.A(sum1[46]), .ZN(n_233));
   INV_X1 i_297 (.A(n_129), .ZN(n_234));
   INV_X1 i_298 (.A(n_125), .ZN(n_235));
   INV_X1 i_299 (.A(sum1[56]), .ZN(n_236));
   INV_X1 i_300 (.A(sum1[57]), .ZN(n_237));
   INV_X1 i_301 (.A(sum1[58]), .ZN(n_238));
   INV_X1 i_302 (.A(sum1[61]), .ZN(n_239));
endmodule

module TreeMultiplierCirc(a, b, out);
   input [31:0]a;
   input [31:0]b;
   output [63:0]out;

   wire [31:0]\c1[1] ;
   wire n_39_0;
   wire n_39_1;
   wire n_39_2;
   wire n_39_3;
   wire n_39_4;
   wire n_39_5;
   wire n_39_6;
   wire n_39_7;
   wire n_39_8;
   wire n_39_9;
   wire n_39_10;
   wire n_39_11;
   wire n_39_12;
   wire n_39_13;
   wire n_39_14;
   wire n_39_15;
   wire n_39_16;
   wire n_39_17;
   wire n_39_18;
   wire n_39_19;
   wire n_39_20;
   wire n_39_21;
   wire n_39_22;
   wire n_39_23;
   wire n_39_24;
   wire n_39_25;
   wire n_39_26;
   wire n_39_27;
   wire n_39_28;
   wire n_39_29;
   wire n_39_30;
   wire [31:0]\c1[2] ;
   wire n_39_32;
   wire n_39_33;
   wire n_39_34;
   wire n_39_35;
   wire n_39_36;
   wire n_39_37;
   wire n_39_38;
   wire n_39_39;
   wire n_39_40;
   wire n_39_41;
   wire n_39_42;
   wire n_39_43;
   wire n_39_44;
   wire n_39_45;
   wire n_39_46;
   wire n_39_47;
   wire n_39_48;
   wire n_39_49;
   wire n_39_50;
   wire n_39_51;
   wire n_39_52;
   wire n_39_53;
   wire n_39_54;
   wire n_39_55;
   wire n_39_56;
   wire n_39_57;
   wire n_39_58;
   wire n_39_59;
   wire n_39_60;
   wire n_39_61;
   wire n_39_62;
   wire [31:0]\c1[3] ;
   wire n_39_64;
   wire n_39_65;
   wire n_39_66;
   wire n_39_67;
   wire n_39_68;
   wire n_39_69;
   wire n_39_70;
   wire n_39_71;
   wire n_39_72;
   wire n_39_73;
   wire n_39_74;
   wire n_39_75;
   wire n_39_76;
   wire n_39_77;
   wire n_39_78;
   wire n_39_79;
   wire n_39_80;
   wire n_39_81;
   wire n_39_82;
   wire n_39_83;
   wire n_39_84;
   wire n_39_85;
   wire n_39_86;
   wire n_39_87;
   wire n_39_88;
   wire n_39_89;
   wire n_39_90;
   wire n_39_91;
   wire n_39_92;
   wire n_39_93;
   wire n_39_94;
   wire [31:0]\c1[4] ;
   wire n_39_96;
   wire n_39_97;
   wire n_39_98;
   wire n_39_99;
   wire n_39_100;
   wire n_39_101;
   wire n_39_102;
   wire n_39_103;
   wire n_39_104;
   wire n_39_105;
   wire n_39_106;
   wire n_39_107;
   wire n_39_108;
   wire n_39_109;
   wire n_39_110;
   wire n_39_111;
   wire n_39_112;
   wire n_39_113;
   wire n_39_114;
   wire n_39_115;
   wire n_39_116;
   wire n_39_117;
   wire n_39_118;
   wire n_39_119;
   wire n_39_120;
   wire n_39_121;
   wire n_39_122;
   wire n_39_123;
   wire n_39_124;
   wire n_39_125;
   wire n_39_126;
   wire [31:0]\c1[5] ;
   wire n_39_128;
   wire n_39_129;
   wire n_39_130;
   wire n_39_131;
   wire n_39_132;
   wire n_39_133;
   wire n_39_134;
   wire n_39_135;
   wire n_39_136;
   wire n_39_137;
   wire n_39_138;
   wire n_39_139;
   wire n_39_140;
   wire n_39_141;
   wire n_39_142;
   wire n_39_143;
   wire n_39_144;
   wire n_39_145;
   wire n_39_146;
   wire n_39_147;
   wire n_39_148;
   wire n_39_149;
   wire n_39_150;
   wire n_39_151;
   wire n_39_152;
   wire n_39_153;
   wire n_39_154;
   wire n_39_155;
   wire n_39_156;
   wire n_39_157;
   wire n_39_158;
   wire [31:0]\c1[6] ;
   wire n_39_160;
   wire n_39_161;
   wire n_39_162;
   wire n_39_163;
   wire n_39_164;
   wire n_39_165;
   wire n_39_166;
   wire n_39_167;
   wire n_39_168;
   wire n_39_169;
   wire n_39_170;
   wire n_39_171;
   wire n_39_172;
   wire n_39_173;
   wire n_39_174;
   wire n_39_175;
   wire n_39_176;
   wire n_39_177;
   wire n_39_178;
   wire n_39_179;
   wire n_39_180;
   wire n_39_181;
   wire n_39_182;
   wire n_39_183;
   wire n_39_184;
   wire n_39_185;
   wire n_39_186;
   wire n_39_187;
   wire n_39_188;
   wire n_39_189;
   wire n_39_190;
   wire [31:0]\c1[7] ;
   wire n_39_192;
   wire n_39_193;
   wire n_39_194;
   wire n_39_195;
   wire n_39_196;
   wire n_39_197;
   wire n_39_198;
   wire n_39_199;
   wire n_39_200;
   wire n_39_201;
   wire n_39_202;
   wire n_39_203;
   wire n_39_204;
   wire n_39_205;
   wire n_39_206;
   wire n_39_207;
   wire n_39_208;
   wire n_39_209;
   wire n_39_210;
   wire n_39_211;
   wire n_39_212;
   wire n_39_213;
   wire n_39_214;
   wire n_39_215;
   wire n_39_216;
   wire n_39_217;
   wire n_39_218;
   wire n_39_219;
   wire n_39_220;
   wire n_39_221;
   wire n_39_222;
   wire [31:0]\c1[8] ;
   wire n_39_224;
   wire n_39_225;
   wire n_39_226;
   wire n_39_227;
   wire n_39_228;
   wire n_39_229;
   wire n_39_230;
   wire n_39_231;
   wire n_39_232;
   wire n_39_233;
   wire n_39_234;
   wire n_39_235;
   wire n_39_236;
   wire n_39_237;
   wire n_39_238;
   wire n_39_239;
   wire n_39_240;
   wire n_39_241;
   wire n_39_242;
   wire n_39_243;
   wire n_39_244;
   wire n_39_245;
   wire n_39_246;
   wire n_39_247;
   wire n_39_248;
   wire n_39_249;
   wire n_39_250;
   wire n_39_251;
   wire n_39_252;
   wire n_39_253;
   wire n_39_254;
   wire [31:0]\c1[9] ;
   wire n_39_256;
   wire n_39_257;
   wire n_39_258;
   wire n_39_259;
   wire n_39_260;
   wire n_39_261;
   wire n_39_262;
   wire n_39_263;
   wire n_39_264;
   wire n_39_265;
   wire n_39_266;
   wire n_39_267;
   wire n_39_268;
   wire n_39_269;
   wire n_39_270;
   wire n_39_271;
   wire n_39_272;
   wire n_39_273;
   wire n_39_274;
   wire n_39_275;
   wire n_39_276;
   wire n_39_277;
   wire n_39_278;
   wire n_39_279;
   wire n_39_280;
   wire n_39_281;
   wire n_39_282;
   wire n_39_283;
   wire n_39_284;
   wire n_39_285;
   wire n_39_286;
   wire [31:0]\c1[10] ;
   wire n_39_288;
   wire n_39_289;
   wire n_39_290;
   wire n_39_291;
   wire n_39_292;
   wire n_39_293;
   wire n_39_294;
   wire n_39_295;
   wire n_39_296;
   wire n_39_297;
   wire n_39_298;
   wire n_39_299;
   wire n_39_300;
   wire n_39_301;
   wire n_39_302;
   wire n_39_303;
   wire n_39_304;
   wire n_39_305;
   wire n_39_306;
   wire n_39_307;
   wire n_39_308;
   wire n_39_309;
   wire n_39_310;
   wire n_39_311;
   wire n_39_312;
   wire n_39_313;
   wire n_39_314;
   wire n_39_315;
   wire n_39_316;
   wire n_39_317;
   wire n_39_318;
   wire [31:0]\c1[11] ;
   wire n_39_320;
   wire n_39_321;
   wire n_39_322;
   wire n_39_323;
   wire n_39_324;
   wire n_39_325;
   wire n_39_326;
   wire n_39_327;
   wire n_39_328;
   wire n_39_329;
   wire n_39_330;
   wire n_39_331;
   wire n_39_332;
   wire n_39_333;
   wire n_39_334;
   wire n_39_335;
   wire n_39_336;
   wire n_39_337;
   wire n_39_338;
   wire n_39_339;
   wire n_39_340;
   wire n_39_341;
   wire n_39_342;
   wire n_39_343;
   wire n_39_344;
   wire n_39_345;
   wire n_39_346;
   wire n_39_347;
   wire n_39_348;
   wire n_39_349;
   wire n_39_350;
   wire [31:0]\c1[12] ;
   wire n_39_352;
   wire n_39_353;
   wire n_39_354;
   wire n_39_355;
   wire n_39_356;
   wire n_39_357;
   wire n_39_358;
   wire n_39_359;
   wire n_39_360;
   wire n_39_361;
   wire n_39_362;
   wire n_39_363;
   wire n_39_364;
   wire n_39_365;
   wire n_39_366;
   wire n_39_367;
   wire n_39_368;
   wire n_39_369;
   wire n_39_370;
   wire n_39_371;
   wire n_39_372;
   wire n_39_373;
   wire n_39_374;
   wire n_39_375;
   wire n_39_376;
   wire n_39_377;
   wire n_39_378;
   wire n_39_379;
   wire n_39_380;
   wire n_39_381;
   wire n_39_382;
   wire [31:0]\c1[13] ;
   wire n_39_384;
   wire n_39_385;
   wire n_39_386;
   wire n_39_387;
   wire n_39_388;
   wire n_39_389;
   wire n_39_390;
   wire n_39_391;
   wire n_39_392;
   wire n_39_393;
   wire n_39_394;
   wire n_39_395;
   wire n_39_396;
   wire n_39_397;
   wire n_39_398;
   wire n_39_399;
   wire n_39_400;
   wire n_39_401;
   wire n_39_402;
   wire n_39_403;
   wire n_39_404;
   wire n_39_405;
   wire n_39_406;
   wire n_39_407;
   wire n_39_408;
   wire n_39_409;
   wire n_39_410;
   wire n_39_411;
   wire n_39_412;
   wire n_39_413;
   wire n_39_414;
   wire [31:0]\c1[14] ;
   wire n_39_416;
   wire n_39_417;
   wire n_39_418;
   wire n_39_419;
   wire n_39_420;
   wire n_39_421;
   wire n_39_422;
   wire n_39_423;
   wire n_39_424;
   wire n_39_425;
   wire n_39_426;
   wire n_39_427;
   wire n_39_428;
   wire n_39_429;
   wire n_39_430;
   wire n_39_431;
   wire n_39_432;
   wire n_39_433;
   wire n_39_434;
   wire n_39_435;
   wire n_39_436;
   wire n_39_437;
   wire n_39_438;
   wire n_39_439;
   wire n_39_440;
   wire n_39_441;
   wire n_39_442;
   wire n_39_443;
   wire n_39_444;
   wire n_39_445;
   wire n_39_446;
   wire [31:0]\c1[15] ;
   wire n_39_448;
   wire n_39_449;
   wire n_39_450;
   wire n_39_451;
   wire n_39_452;
   wire n_39_453;
   wire n_39_454;
   wire n_39_455;
   wire n_39_456;
   wire n_39_457;
   wire n_39_458;
   wire n_39_459;
   wire n_39_460;
   wire n_39_461;
   wire n_39_462;
   wire n_39_463;
   wire n_39_464;
   wire n_39_465;
   wire n_39_466;
   wire n_39_467;
   wire n_39_468;
   wire n_39_469;
   wire n_39_470;
   wire n_39_471;
   wire n_39_472;
   wire n_39_473;
   wire n_39_474;
   wire n_39_475;
   wire n_39_476;
   wire n_39_477;
   wire n_39_478;
   wire [31:0]\c1[16] ;
   wire n_39_480;
   wire n_39_481;
   wire n_39_482;
   wire n_39_483;
   wire n_39_484;
   wire n_39_485;
   wire n_39_486;
   wire n_39_487;
   wire n_39_488;
   wire n_39_489;
   wire n_39_490;
   wire n_39_491;
   wire n_39_492;
   wire n_39_493;
   wire n_39_494;
   wire n_39_495;
   wire n_39_496;
   wire n_39_497;
   wire n_39_498;
   wire n_39_499;
   wire n_39_500;
   wire n_39_501;
   wire n_39_502;
   wire n_39_503;
   wire n_39_504;
   wire n_39_505;
   wire n_39_506;
   wire n_39_507;
   wire n_39_508;
   wire n_39_509;
   wire n_39_510;
   wire [31:0]\c1[17] ;
   wire n_39_512;
   wire n_39_513;
   wire n_39_514;
   wire n_39_515;
   wire n_39_516;
   wire n_39_517;
   wire n_39_518;
   wire n_39_519;
   wire n_39_520;
   wire n_39_521;
   wire n_39_522;
   wire n_39_523;
   wire n_39_524;
   wire n_39_525;
   wire n_39_526;
   wire n_39_527;
   wire n_39_528;
   wire n_39_529;
   wire n_39_530;
   wire n_39_531;
   wire n_39_532;
   wire n_39_533;
   wire n_39_534;
   wire n_39_535;
   wire n_39_536;
   wire n_39_537;
   wire n_39_538;
   wire n_39_539;
   wire n_39_540;
   wire n_39_541;
   wire n_39_542;
   wire [31:0]\c1[18] ;
   wire n_39_544;
   wire n_39_545;
   wire n_39_546;
   wire n_39_547;
   wire n_39_548;
   wire n_39_549;
   wire n_39_550;
   wire n_39_551;
   wire n_39_552;
   wire n_39_553;
   wire n_39_554;
   wire n_39_555;
   wire n_39_556;
   wire n_39_557;
   wire n_39_558;
   wire n_39_559;
   wire n_39_560;
   wire n_39_561;
   wire n_39_562;
   wire n_39_563;
   wire n_39_564;
   wire n_39_565;
   wire n_39_566;
   wire n_39_567;
   wire n_39_568;
   wire n_39_569;
   wire n_39_570;
   wire n_39_571;
   wire n_39_572;
   wire n_39_573;
   wire n_39_574;
   wire [31:0]\c1[19] ;
   wire n_39_576;
   wire n_39_577;
   wire n_39_578;
   wire n_39_579;
   wire n_39_580;
   wire n_39_581;
   wire n_39_582;
   wire n_39_583;
   wire n_39_584;
   wire n_39_585;
   wire n_39_586;
   wire n_39_587;
   wire n_39_588;
   wire n_39_589;
   wire n_39_590;
   wire n_39_591;
   wire n_39_592;
   wire n_39_593;
   wire n_39_594;
   wire n_39_595;
   wire n_39_596;
   wire n_39_597;
   wire n_39_598;
   wire n_39_599;
   wire n_39_600;
   wire n_39_601;
   wire n_39_602;
   wire n_39_603;
   wire n_39_604;
   wire n_39_605;
   wire n_39_606;
   wire [31:0]\c1[20] ;
   wire n_39_608;
   wire n_39_609;
   wire n_39_610;
   wire n_39_611;
   wire n_39_612;
   wire n_39_613;
   wire n_39_614;
   wire n_39_615;
   wire n_39_616;
   wire n_39_617;
   wire n_39_618;
   wire n_39_619;
   wire n_39_620;
   wire n_39_621;
   wire n_39_622;
   wire n_39_623;
   wire n_39_624;
   wire n_39_625;
   wire n_39_626;
   wire n_39_627;
   wire n_39_628;
   wire n_39_629;
   wire n_39_630;
   wire n_39_631;
   wire n_39_632;
   wire n_39_633;
   wire n_39_634;
   wire n_39_635;
   wire n_39_636;
   wire n_39_637;
   wire n_39_638;
   wire [31:0]\c1[21] ;
   wire n_39_640;
   wire n_39_641;
   wire n_39_642;
   wire n_39_643;
   wire n_39_644;
   wire n_39_645;
   wire n_39_646;
   wire n_39_647;
   wire n_39_648;
   wire n_39_649;
   wire n_39_650;
   wire n_39_651;
   wire n_39_652;
   wire n_39_653;
   wire n_39_654;
   wire n_39_655;
   wire n_39_656;
   wire n_39_657;
   wire n_39_658;
   wire n_39_659;
   wire n_39_660;
   wire n_39_661;
   wire n_39_662;
   wire n_39_663;
   wire n_39_664;
   wire n_39_665;
   wire n_39_666;
   wire n_39_667;
   wire n_39_668;
   wire n_39_669;
   wire n_39_670;
   wire [31:0]\c1[22] ;
   wire n_39_672;
   wire n_39_673;
   wire n_39_674;
   wire n_39_675;
   wire n_39_676;
   wire n_39_677;
   wire n_39_678;
   wire n_39_679;
   wire n_39_680;
   wire n_39_681;
   wire n_39_682;
   wire n_39_683;
   wire n_39_684;
   wire n_39_685;
   wire n_39_686;
   wire n_39_687;
   wire n_39_688;
   wire n_39_689;
   wire n_39_690;
   wire n_39_691;
   wire n_39_692;
   wire n_39_693;
   wire n_39_694;
   wire n_39_695;
   wire n_39_696;
   wire n_39_697;
   wire n_39_698;
   wire n_39_699;
   wire n_39_700;
   wire n_39_701;
   wire n_39_702;
   wire [31:0]\c1[23] ;
   wire n_39_704;
   wire n_39_705;
   wire n_39_706;
   wire n_39_707;
   wire n_39_708;
   wire n_39_709;
   wire n_39_710;
   wire n_39_711;
   wire n_39_712;
   wire n_39_713;
   wire n_39_714;
   wire n_39_715;
   wire n_39_716;
   wire n_39_717;
   wire n_39_718;
   wire n_39_719;
   wire n_39_720;
   wire n_39_721;
   wire n_39_722;
   wire n_39_723;
   wire n_39_724;
   wire n_39_725;
   wire n_39_726;
   wire n_39_727;
   wire n_39_728;
   wire n_39_729;
   wire n_39_730;
   wire n_39_731;
   wire n_39_732;
   wire n_39_733;
   wire n_39_734;
   wire [31:0]\c1[24] ;
   wire n_39_736;
   wire n_39_737;
   wire n_39_738;
   wire n_39_739;
   wire n_39_740;
   wire n_39_741;
   wire n_39_742;
   wire n_39_743;
   wire n_39_744;
   wire n_39_745;
   wire n_39_746;
   wire n_39_747;
   wire n_39_748;
   wire n_39_749;
   wire n_39_750;
   wire n_39_751;
   wire n_39_752;
   wire n_39_753;
   wire n_39_754;
   wire n_39_755;
   wire n_39_756;
   wire n_39_757;
   wire n_39_758;
   wire n_39_759;
   wire n_39_760;
   wire n_39_761;
   wire n_39_762;
   wire n_39_763;
   wire n_39_764;
   wire n_39_765;
   wire n_39_766;
   wire [31:0]\c1[25] ;
   wire n_39_768;
   wire n_39_769;
   wire n_39_770;
   wire n_39_771;
   wire n_39_772;
   wire n_39_773;
   wire n_39_774;
   wire n_39_775;
   wire n_39_776;
   wire n_39_777;
   wire n_39_778;
   wire n_39_779;
   wire n_39_780;
   wire n_39_781;
   wire n_39_782;
   wire n_39_783;
   wire n_39_784;
   wire n_39_785;
   wire n_39_786;
   wire n_39_787;
   wire n_39_788;
   wire n_39_789;
   wire n_39_790;
   wire n_39_791;
   wire n_39_792;
   wire n_39_793;
   wire n_39_794;
   wire n_39_795;
   wire n_39_796;
   wire n_39_797;
   wire n_39_798;
   wire [31:0]\c1[26] ;
   wire n_39_800;
   wire n_39_801;
   wire n_39_802;
   wire n_39_803;
   wire n_39_804;
   wire n_39_805;
   wire n_39_806;
   wire n_39_807;
   wire n_39_808;
   wire n_39_809;
   wire n_39_810;
   wire n_39_811;
   wire n_39_812;
   wire n_39_813;
   wire n_39_814;
   wire n_39_815;
   wire n_39_816;
   wire n_39_817;
   wire n_39_818;
   wire n_39_819;
   wire n_39_820;
   wire n_39_821;
   wire n_39_822;
   wire n_39_823;
   wire n_39_824;
   wire n_39_825;
   wire n_39_826;
   wire n_39_827;
   wire n_39_828;
   wire n_39_829;
   wire n_39_830;
   wire [31:0]\c1[27] ;
   wire n_39_832;
   wire n_39_833;
   wire n_39_834;
   wire n_39_835;
   wire n_39_836;
   wire n_39_837;
   wire n_39_838;
   wire n_39_839;
   wire n_39_840;
   wire n_39_841;
   wire n_39_842;
   wire n_39_843;
   wire n_39_844;
   wire n_39_845;
   wire n_39_846;
   wire n_39_847;
   wire n_39_848;
   wire n_39_849;
   wire n_39_850;
   wire n_39_851;
   wire n_39_852;
   wire n_39_853;
   wire n_39_854;
   wire n_39_855;
   wire n_39_856;
   wire n_39_857;
   wire n_39_858;
   wire n_39_859;
   wire n_39_860;
   wire n_39_861;
   wire n_39_862;
   wire [31:0]\c1[28] ;
   wire n_39_864;
   wire n_39_865;
   wire n_39_866;
   wire n_39_867;
   wire n_39_31;
   wire n_39_63;
   wire n_39_95;
   wire n_39_127;
   wire n_39_159;
   wire n_39_191;
   wire n_39_223;
   wire n_39_255;
   wire n_39_287;
   wire n_39_319;
   wire n_39_351;
   wire n_39_383;
   wire n_39_415;
   wire n_39_447;
   wire n_39_479;
   wire n_39_511;
   wire n_39_543;
   wire n_39_575;
   wire n_39_607;
   wire n_39_639;
   wire n_39_671;
   wire n_39_703;
   wire n_39_735;
   wire n_39_767;
   wire n_39_799;
   wire n_39_831;
   wire n_39_863;
   wire [31:0]\c1[29] ;
   wire [32:0]\s1[29] ;
   wire n_4_0_1;
   wire n_4_0_2;
   wire [31:0]\partial_reg[0] ;
   wire n_4_0_3;
   wire n_4_0_4;
   wire n_4_0_5;
   wire n_4_0_6;
   wire n_4_0_7;
   wire n_4_0_8;
   wire n_4_0_9;
   wire n_4_0_10;
   wire n_4_0_11;
   wire n_4_0_12;
   wire n_4_0_13;
   wire n_4_0_14;
   wire n_4_0_15;
   wire n_4_0_16;
   wire n_4_0_17;
   wire n_4_0_18;
   wire n_4_0_19;
   wire n_4_0_20;
   wire n_4_0_21;
   wire n_4_0_22;
   wire n_4_0_23;
   wire n_4_0_24;
   wire n_4_0_25;
   wire n_4_0_26;
   wire n_4_0_27;
   wire n_4_0_28;
   wire n_4_0_29;
   wire [31:0]\partial_reg[1] ;
   wire [31:0]\partial_reg[2] ;
   wire n_4_0_35;
   wire [31:0]\partial_reg[3] ;
   wire n_4_0_36;
   wire [31:0]\partial_reg[4] ;
   wire n_4_0_37;
   wire [31:0]\partial_reg[5] ;
   wire n_4_0_38;
   wire [31:0]\partial_reg[6] ;
   wire n_4_0_39;
   wire [31:0]\partial_reg[7] ;
   wire n_4_0_40;
   wire [31:0]\partial_reg[8] ;
   wire n_4_0_41;
   wire [31:0]\partial_reg[9] ;
   wire n_4_0_42;
   wire [31:0]\partial_reg[10] ;
   wire n_4_0_43;
   wire [31:0]\partial_reg[11] ;
   wire n_4_0_44;
   wire [31:0]\partial_reg[12] ;
   wire n_4_0_45;
   wire [31:0]\partial_reg[13] ;
   wire n_4_0_46;
   wire [31:0]\partial_reg[14] ;
   wire n_4_0_47;
   wire [31:0]\partial_reg[15] ;
   wire n_4_0_48;
   wire [31:0]\partial_reg[16] ;
   wire n_4_0_49;
   wire [31:0]\partial_reg[17] ;
   wire n_4_0_50;
   wire [31:0]\partial_reg[18] ;
   wire n_4_0_51;
   wire [31:0]\partial_reg[19] ;
   wire n_4_0_52;
   wire [31:0]\partial_reg[20] ;
   wire n_4_0_53;
   wire [31:0]\partial_reg[21] ;
   wire n_4_0_54;
   wire [31:0]\partial_reg[22] ;
   wire n_4_0_55;
   wire [31:0]\partial_reg[23] ;
   wire n_4_0_56;
   wire [31:0]\partial_reg[24] ;
   wire n_4_0_57;
   wire [31:0]\partial_reg[25] ;
   wire n_4_0_58;
   wire [31:0]\partial_reg[26] ;
   wire n_4_0_59;
   wire [31:0]\partial_reg[27] ;
   wire n_4_0_60;
   wire [31:0]\partial_reg[28] ;
   wire n_4_0_61;
   wire [31:0]\partial_reg[29] ;
   wire n_4_0_62;
   wire [31:0]\partial_reg[30] ;
   wire n_4_0_63;
   wire [31:0]\partial_reg[31] ;
   wire n_4_0_34;
   wire n_4_0_33;
   wire n_4_0_32;
   wire n_4_0_31;
   wire n_4_0_30;
   wire n_4_0_0;
   wire n_4_0_64;
   wire n_4_0_65;
   wire [31:0]\c1[0] ;
   wire [32:0]\s1[0] ;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire [31:0]op2;
   wire [31:0]op1;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_1_18;
   wire n_0_1_19;
   wire n_0_1_20;
   wire n_0_1_21;
   wire n_0_1_22;
   wire n_0_1_23;
   wire n_0_1_24;
   wire n_0_1_25;
   wire n_0_1_26;
   wire n_0_1_27;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_1_30;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_11;

   PartialAdder__1_186 genblk1_1_p2 (.a({\partial_reg[2] [31], \s1[0] [31], 
      \s1[0] [30], \s1[0] [29], \s1[0] [28], \s1[0] [27], \s1[0] [26], 
      \s1[0] [25], \s1[0] [24], \s1[0] [23], \s1[0] [22], \s1[0] [21], 
      \s1[0] [20], \s1[0] [19], \s1[0] [18], \s1[0] [17], \s1[0] [16], 
      \s1[0] [15], \s1[0] [14], \s1[0] [13], \s1[0] [12], \s1[0] [11], 
      \s1[0] [10], \s1[0] [9], \s1[0] [8], \s1[0] [7], \s1[0] [6], \s1[0] [5], 
      \s1[0] [4], \s1[0] [3], \s1[0] [2], \s1[0] [1], uc_0}), .b(\c1[0] ), 
      .c({uc_1, \partial_reg[3] [30], \partial_reg[3] [29], \partial_reg[3] [28], 
      \partial_reg[3] [27], \partial_reg[3] [26], \partial_reg[3] [25], 
      \partial_reg[3] [24], \partial_reg[3] [23], \partial_reg[3] [22], 
      \partial_reg[3] [21], \partial_reg[3] [20], \partial_reg[3] [19], 
      \partial_reg[3] [18], \partial_reg[3] [17], \partial_reg[3] [16], 
      \partial_reg[3] [15], \partial_reg[3] [14], \partial_reg[3] [13], 
      \partial_reg[3] [12], \partial_reg[3] [11], \partial_reg[3] [10], 
      \partial_reg[3] [9], \partial_reg[3] [8], \partial_reg[3] [7], 
      \partial_reg[3] [6], \partial_reg[3] [5], \partial_reg[3] [4], 
      \partial_reg[3] [3], \partial_reg[3] [2], \partial_reg[3] [1], 
      \partial_reg[3] [0]}), .s1({uc_2, n_39_30, n_39_29, n_39_28, n_39_27, 
      n_39_26, n_39_25, n_39_24, n_39_23, n_39_22, n_39_21, n_39_20, n_39_19, 
      n_39_18, n_39_17, n_39_16, n_39_15, n_39_14, n_39_13, n_39_12, n_39_11, 
      n_39_10, n_39_9, n_39_8, n_39_7, n_39_6, n_39_5, n_39_4, n_39_3, n_39_2, 
      n_39_1, n_39_0, n_0}), .c1(\c1[1] ));
   PartialAdder__1_283 genblk1_2_p2 (.a({\partial_reg[3] [31], n_39_30, n_39_29, 
      n_39_28, n_39_27, n_39_26, n_39_25, n_39_24, n_39_23, n_39_22, n_39_21, 
      n_39_20, n_39_19, n_39_18, n_39_17, n_39_16, n_39_15, n_39_14, n_39_13, 
      n_39_12, n_39_11, n_39_10, n_39_9, n_39_8, n_39_7, n_39_6, n_39_5, n_39_4, 
      n_39_3, n_39_2, n_39_1, n_39_0, uc_3}), .b(\c1[1] ), .c({uc_4, 
      \partial_reg[4] [30], \partial_reg[4] [29], \partial_reg[4] [28], 
      \partial_reg[4] [27], \partial_reg[4] [26], \partial_reg[4] [25], 
      \partial_reg[4] [24], \partial_reg[4] [23], \partial_reg[4] [22], 
      \partial_reg[4] [21], \partial_reg[4] [20], \partial_reg[4] [19], 
      \partial_reg[4] [18], \partial_reg[4] [17], \partial_reg[4] [16], 
      \partial_reg[4] [15], \partial_reg[4] [14], \partial_reg[4] [13], 
      \partial_reg[4] [12], \partial_reg[4] [11], \partial_reg[4] [10], 
      \partial_reg[4] [9], \partial_reg[4] [8], \partial_reg[4] [7], 
      \partial_reg[4] [6], \partial_reg[4] [5], \partial_reg[4] [4], 
      \partial_reg[4] [3], \partial_reg[4] [2], \partial_reg[4] [1], 
      \partial_reg[4] [0]}), .s1({uc_5, n_39_62, n_39_61, n_39_60, n_39_59, 
      n_39_58, n_39_57, n_39_56, n_39_55, n_39_54, n_39_53, n_39_52, n_39_51, 
      n_39_50, n_39_49, n_39_48, n_39_47, n_39_46, n_39_45, n_39_44, n_39_43, 
      n_39_42, n_39_41, n_39_40, n_39_39, n_39_38, n_39_37, n_39_36, n_39_35, 
      n_39_34, n_39_33, n_39_32, n_1}), .c1(\c1[2] ));
   PartialAdder__1_380 genblk1_3_p2 (.a({\partial_reg[4] [31], n_39_62, n_39_61, 
      n_39_60, n_39_59, n_39_58, n_39_57, n_39_56, n_39_55, n_39_54, n_39_53, 
      n_39_52, n_39_51, n_39_50, n_39_49, n_39_48, n_39_47, n_39_46, n_39_45, 
      n_39_44, n_39_43, n_39_42, n_39_41, n_39_40, n_39_39, n_39_38, n_39_37, 
      n_39_36, n_39_35, n_39_34, n_39_33, n_39_32, uc_6}), .b(\c1[2] ), .c({uc_7, 
      \partial_reg[5] [30], \partial_reg[5] [29], \partial_reg[5] [28], 
      \partial_reg[5] [27], \partial_reg[5] [26], \partial_reg[5] [25], 
      \partial_reg[5] [24], \partial_reg[5] [23], \partial_reg[5] [22], 
      \partial_reg[5] [21], \partial_reg[5] [20], \partial_reg[5] [19], 
      \partial_reg[5] [18], \partial_reg[5] [17], \partial_reg[5] [16], 
      \partial_reg[5] [15], \partial_reg[5] [14], \partial_reg[5] [13], 
      \partial_reg[5] [12], \partial_reg[5] [11], \partial_reg[5] [10], 
      \partial_reg[5] [9], \partial_reg[5] [8], \partial_reg[5] [7], 
      \partial_reg[5] [6], \partial_reg[5] [5], \partial_reg[5] [4], 
      \partial_reg[5] [3], \partial_reg[5] [2], \partial_reg[5] [1], 
      \partial_reg[5] [0]}), .s1({uc_8, n_39_94, n_39_93, n_39_92, n_39_91, 
      n_39_90, n_39_89, n_39_88, n_39_87, n_39_86, n_39_85, n_39_84, n_39_83, 
      n_39_82, n_39_81, n_39_80, n_39_79, n_39_78, n_39_77, n_39_76, n_39_75, 
      n_39_74, n_39_73, n_39_72, n_39_71, n_39_70, n_39_69, n_39_68, n_39_67, 
      n_39_66, n_39_65, n_39_64, n_2}), .c1(\c1[3] ));
   PartialAdder__1_477 genblk1_4_p2 (.a({\partial_reg[5] [31], n_39_94, n_39_93, 
      n_39_92, n_39_91, n_39_90, n_39_89, n_39_88, n_39_87, n_39_86, n_39_85, 
      n_39_84, n_39_83, n_39_82, n_39_81, n_39_80, n_39_79, n_39_78, n_39_77, 
      n_39_76, n_39_75, n_39_74, n_39_73, n_39_72, n_39_71, n_39_70, n_39_69, 
      n_39_68, n_39_67, n_39_66, n_39_65, n_39_64, uc_9}), .b(\c1[3] ), .c({
      uc_10, \partial_reg[6] [30], \partial_reg[6] [29], \partial_reg[6] [28], 
      \partial_reg[6] [27], \partial_reg[6] [26], \partial_reg[6] [25], 
      \partial_reg[6] [24], \partial_reg[6] [23], \partial_reg[6] [22], 
      \partial_reg[6] [21], \partial_reg[6] [20], \partial_reg[6] [19], 
      \partial_reg[6] [18], \partial_reg[6] [17], \partial_reg[6] [16], 
      \partial_reg[6] [15], \partial_reg[6] [14], \partial_reg[6] [13], 
      \partial_reg[6] [12], \partial_reg[6] [11], \partial_reg[6] [10], 
      \partial_reg[6] [9], \partial_reg[6] [8], \partial_reg[6] [7], 
      \partial_reg[6] [6], \partial_reg[6] [5], \partial_reg[6] [4], 
      \partial_reg[6] [3], \partial_reg[6] [2], \partial_reg[6] [1], 
      \partial_reg[6] [0]}), .s1({uc_11, n_39_126, n_39_125, n_39_124, n_39_123, 
      n_39_122, n_39_121, n_39_120, n_39_119, n_39_118, n_39_117, n_39_116, 
      n_39_115, n_39_114, n_39_113, n_39_112, n_39_111, n_39_110, n_39_109, 
      n_39_108, n_39_107, n_39_106, n_39_105, n_39_104, n_39_103, n_39_102, 
      n_39_101, n_39_100, n_39_99, n_39_98, n_39_97, n_39_96, n_3}), .c1(\c1[4] ));
   PartialAdder__1_574 genblk1_5_p2 (.a({\partial_reg[6] [31], n_39_126, 
      n_39_125, n_39_124, n_39_123, n_39_122, n_39_121, n_39_120, n_39_119, 
      n_39_118, n_39_117, n_39_116, n_39_115, n_39_114, n_39_113, n_39_112, 
      n_39_111, n_39_110, n_39_109, n_39_108, n_39_107, n_39_106, n_39_105, 
      n_39_104, n_39_103, n_39_102, n_39_101, n_39_100, n_39_99, n_39_98, 
      n_39_97, n_39_96, uc_12}), .b(\c1[4] ), .c({uc_13, \partial_reg[7] [30], 
      \partial_reg[7] [29], \partial_reg[7] [28], \partial_reg[7] [27], 
      \partial_reg[7] [26], \partial_reg[7] [25], \partial_reg[7] [24], 
      \partial_reg[7] [23], \partial_reg[7] [22], \partial_reg[7] [21], 
      \partial_reg[7] [20], \partial_reg[7] [19], \partial_reg[7] [18], 
      \partial_reg[7] [17], \partial_reg[7] [16], \partial_reg[7] [15], 
      \partial_reg[7] [14], \partial_reg[7] [13], \partial_reg[7] [12], 
      \partial_reg[7] [11], \partial_reg[7] [10], \partial_reg[7] [9], 
      \partial_reg[7] [8], \partial_reg[7] [7], \partial_reg[7] [6], 
      \partial_reg[7] [5], \partial_reg[7] [4], \partial_reg[7] [3], 
      \partial_reg[7] [2], \partial_reg[7] [1], \partial_reg[7] [0]}), .s1({
      uc_14, n_39_158, n_39_157, n_39_156, n_39_155, n_39_154, n_39_153, 
      n_39_152, n_39_151, n_39_150, n_39_149, n_39_148, n_39_147, n_39_146, 
      n_39_145, n_39_144, n_39_143, n_39_142, n_39_141, n_39_140, n_39_139, 
      n_39_138, n_39_137, n_39_136, n_39_135, n_39_134, n_39_133, n_39_132, 
      n_39_131, n_39_130, n_39_129, n_39_128, n_4}), .c1(\c1[5] ));
   PartialAdder__1_671 genblk1_6_p2 (.a({\partial_reg[7] [31], n_39_158, 
      n_39_157, n_39_156, n_39_155, n_39_154, n_39_153, n_39_152, n_39_151, 
      n_39_150, n_39_149, n_39_148, n_39_147, n_39_146, n_39_145, n_39_144, 
      n_39_143, n_39_142, n_39_141, n_39_140, n_39_139, n_39_138, n_39_137, 
      n_39_136, n_39_135, n_39_134, n_39_133, n_39_132, n_39_131, n_39_130, 
      n_39_129, n_39_128, uc_15}), .b(\c1[5] ), .c({uc_16, \partial_reg[8] [30], 
      \partial_reg[8] [29], \partial_reg[8] [28], \partial_reg[8] [27], 
      \partial_reg[8] [26], \partial_reg[8] [25], \partial_reg[8] [24], 
      \partial_reg[8] [23], \partial_reg[8] [22], \partial_reg[8] [21], 
      \partial_reg[8] [20], \partial_reg[8] [19], \partial_reg[8] [18], 
      \partial_reg[8] [17], \partial_reg[8] [16], \partial_reg[8] [15], 
      \partial_reg[8] [14], \partial_reg[8] [13], \partial_reg[8] [12], 
      \partial_reg[8] [11], \partial_reg[8] [10], \partial_reg[8] [9], 
      \partial_reg[8] [8], \partial_reg[8] [7], \partial_reg[8] [6], 
      \partial_reg[8] [5], \partial_reg[8] [4], \partial_reg[8] [3], 
      \partial_reg[8] [2], \partial_reg[8] [1], \partial_reg[8] [0]}), .s1({
      uc_17, n_39_190, n_39_189, n_39_188, n_39_187, n_39_186, n_39_185, 
      n_39_184, n_39_183, n_39_182, n_39_181, n_39_180, n_39_179, n_39_178, 
      n_39_177, n_39_176, n_39_175, n_39_174, n_39_173, n_39_172, n_39_171, 
      n_39_170, n_39_169, n_39_168, n_39_167, n_39_166, n_39_165, n_39_164, 
      n_39_163, n_39_162, n_39_161, n_39_160, n_5}), .c1(\c1[6] ));
   PartialAdder__1_768 genblk1_7_p2 (.a({\partial_reg[8] [31], n_39_190, 
      n_39_189, n_39_188, n_39_187, n_39_186, n_39_185, n_39_184, n_39_183, 
      n_39_182, n_39_181, n_39_180, n_39_179, n_39_178, n_39_177, n_39_176, 
      n_39_175, n_39_174, n_39_173, n_39_172, n_39_171, n_39_170, n_39_169, 
      n_39_168, n_39_167, n_39_166, n_39_165, n_39_164, n_39_163, n_39_162, 
      n_39_161, n_39_160, uc_18}), .b(\c1[6] ), .c({uc_19, \partial_reg[9] [30], 
      \partial_reg[9] [29], \partial_reg[9] [28], \partial_reg[9] [27], 
      \partial_reg[9] [26], \partial_reg[9] [25], \partial_reg[9] [24], 
      \partial_reg[9] [23], \partial_reg[9] [22], \partial_reg[9] [21], 
      \partial_reg[9] [20], \partial_reg[9] [19], \partial_reg[9] [18], 
      \partial_reg[9] [17], \partial_reg[9] [16], \partial_reg[9] [15], 
      \partial_reg[9] [14], \partial_reg[9] [13], \partial_reg[9] [12], 
      \partial_reg[9] [11], \partial_reg[9] [10], \partial_reg[9] [9], 
      \partial_reg[9] [8], \partial_reg[9] [7], \partial_reg[9] [6], 
      \partial_reg[9] [5], \partial_reg[9] [4], \partial_reg[9] [3], 
      \partial_reg[9] [2], \partial_reg[9] [1], \partial_reg[9] [0]}), .s1({
      uc_20, n_39_222, n_39_221, n_39_220, n_39_219, n_39_218, n_39_217, 
      n_39_216, n_39_215, n_39_214, n_39_213, n_39_212, n_39_211, n_39_210, 
      n_39_209, n_39_208, n_39_207, n_39_206, n_39_205, n_39_204, n_39_203, 
      n_39_202, n_39_201, n_39_200, n_39_199, n_39_198, n_39_197, n_39_196, 
      n_39_195, n_39_194, n_39_193, n_39_192, n_6}), .c1(\c1[7] ));
   PartialAdder__1_865 genblk1_8_p2 (.a({\partial_reg[9] [31], n_39_222, 
      n_39_221, n_39_220, n_39_219, n_39_218, n_39_217, n_39_216, n_39_215, 
      n_39_214, n_39_213, n_39_212, n_39_211, n_39_210, n_39_209, n_39_208, 
      n_39_207, n_39_206, n_39_205, n_39_204, n_39_203, n_39_202, n_39_201, 
      n_39_200, n_39_199, n_39_198, n_39_197, n_39_196, n_39_195, n_39_194, 
      n_39_193, n_39_192, uc_21}), .b(\c1[7] ), .c({uc_22, \partial_reg[10] [30], 
      \partial_reg[10] [29], \partial_reg[10] [28], \partial_reg[10] [27], 
      \partial_reg[10] [26], \partial_reg[10] [25], \partial_reg[10] [24], 
      \partial_reg[10] [23], \partial_reg[10] [22], \partial_reg[10] [21], 
      \partial_reg[10] [20], \partial_reg[10] [19], \partial_reg[10] [18], 
      \partial_reg[10] [17], \partial_reg[10] [16], \partial_reg[10] [15], 
      \partial_reg[10] [14], \partial_reg[10] [13], \partial_reg[10] [12], 
      \partial_reg[10] [11], \partial_reg[10] [10], \partial_reg[10] [9], 
      \partial_reg[10] [8], \partial_reg[10] [7], \partial_reg[10] [6], 
      \partial_reg[10] [5], \partial_reg[10] [4], \partial_reg[10] [3], 
      \partial_reg[10] [2], \partial_reg[10] [1], \partial_reg[10] [0]}), 
      .s1({uc_23, n_39_254, n_39_253, n_39_252, n_39_251, n_39_250, n_39_249, 
      n_39_248, n_39_247, n_39_246, n_39_245, n_39_244, n_39_243, n_39_242, 
      n_39_241, n_39_240, n_39_239, n_39_238, n_39_237, n_39_236, n_39_235, 
      n_39_234, n_39_233, n_39_232, n_39_231, n_39_230, n_39_229, n_39_228, 
      n_39_227, n_39_226, n_39_225, n_39_224, n_7}), .c1(\c1[8] ));
   PartialAdder__1_962 genblk1_9_p2 (.a({\partial_reg[10] [31], n_39_254, 
      n_39_253, n_39_252, n_39_251, n_39_250, n_39_249, n_39_248, n_39_247, 
      n_39_246, n_39_245, n_39_244, n_39_243, n_39_242, n_39_241, n_39_240, 
      n_39_239, n_39_238, n_39_237, n_39_236, n_39_235, n_39_234, n_39_233, 
      n_39_232, n_39_231, n_39_230, n_39_229, n_39_228, n_39_227, n_39_226, 
      n_39_225, n_39_224, uc_24}), .b(\c1[8] ), .c({uc_25, \partial_reg[11] [30], 
      \partial_reg[11] [29], \partial_reg[11] [28], \partial_reg[11] [27], 
      \partial_reg[11] [26], \partial_reg[11] [25], \partial_reg[11] [24], 
      \partial_reg[11] [23], \partial_reg[11] [22], \partial_reg[11] [21], 
      \partial_reg[11] [20], \partial_reg[11] [19], \partial_reg[11] [18], 
      \partial_reg[11] [17], \partial_reg[11] [16], \partial_reg[11] [15], 
      \partial_reg[11] [14], \partial_reg[11] [13], \partial_reg[11] [12], 
      \partial_reg[11] [11], \partial_reg[11] [10], \partial_reg[11] [9], 
      \partial_reg[11] [8], \partial_reg[11] [7], \partial_reg[11] [6], 
      \partial_reg[11] [5], \partial_reg[11] [4], \partial_reg[11] [3], 
      \partial_reg[11] [2], \partial_reg[11] [1], \partial_reg[11] [0]}), 
      .s1({uc_26, n_39_286, n_39_285, n_39_284, n_39_283, n_39_282, n_39_281, 
      n_39_280, n_39_279, n_39_278, n_39_277, n_39_276, n_39_275, n_39_274, 
      n_39_273, n_39_272, n_39_271, n_39_270, n_39_269, n_39_268, n_39_267, 
      n_39_266, n_39_265, n_39_264, n_39_263, n_39_262, n_39_261, n_39_260, 
      n_39_259, n_39_258, n_39_257, n_39_256, n_8}), .c1(\c1[9] ));
   PartialAdder__1_1059 genblk1_10_p2 (.a({\partial_reg[11] [31], n_39_286, 
      n_39_285, n_39_284, n_39_283, n_39_282, n_39_281, n_39_280, n_39_279, 
      n_39_278, n_39_277, n_39_276, n_39_275, n_39_274, n_39_273, n_39_272, 
      n_39_271, n_39_270, n_39_269, n_39_268, n_39_267, n_39_266, n_39_265, 
      n_39_264, n_39_263, n_39_262, n_39_261, n_39_260, n_39_259, n_39_258, 
      n_39_257, n_39_256, uc_27}), .b(\c1[9] ), .c({uc_28, \partial_reg[12] [30], 
      \partial_reg[12] [29], \partial_reg[12] [28], \partial_reg[12] [27], 
      \partial_reg[12] [26], \partial_reg[12] [25], \partial_reg[12] [24], 
      \partial_reg[12] [23], \partial_reg[12] [22], \partial_reg[12] [21], 
      \partial_reg[12] [20], \partial_reg[12] [19], \partial_reg[12] [18], 
      \partial_reg[12] [17], \partial_reg[12] [16], \partial_reg[12] [15], 
      \partial_reg[12] [14], \partial_reg[12] [13], \partial_reg[12] [12], 
      \partial_reg[12] [11], \partial_reg[12] [10], \partial_reg[12] [9], 
      \partial_reg[12] [8], \partial_reg[12] [7], \partial_reg[12] [6], 
      \partial_reg[12] [5], \partial_reg[12] [4], \partial_reg[12] [3], 
      \partial_reg[12] [2], \partial_reg[12] [1], \partial_reg[12] [0]}), 
      .s1({uc_29, n_39_318, n_39_317, n_39_316, n_39_315, n_39_314, n_39_313, 
      n_39_312, n_39_311, n_39_310, n_39_309, n_39_308, n_39_307, n_39_306, 
      n_39_305, n_39_304, n_39_303, n_39_302, n_39_301, n_39_300, n_39_299, 
      n_39_298, n_39_297, n_39_296, n_39_295, n_39_294, n_39_293, n_39_292, 
      n_39_291, n_39_290, n_39_289, n_39_288, n_9}), .c1(\c1[10] ));
   PartialAdder__1_1156 genblk1_11_p2 (.a({\partial_reg[12] [31], n_39_318, 
      n_39_317, n_39_316, n_39_315, n_39_314, n_39_313, n_39_312, n_39_311, 
      n_39_310, n_39_309, n_39_308, n_39_307, n_39_306, n_39_305, n_39_304, 
      n_39_303, n_39_302, n_39_301, n_39_300, n_39_299, n_39_298, n_39_297, 
      n_39_296, n_39_295, n_39_294, n_39_293, n_39_292, n_39_291, n_39_290, 
      n_39_289, n_39_288, uc_30}), .b(\c1[10] ), .c({uc_31, 
      \partial_reg[13] [30], \partial_reg[13] [29], \partial_reg[13] [28], 
      \partial_reg[13] [27], \partial_reg[13] [26], \partial_reg[13] [25], 
      \partial_reg[13] [24], \partial_reg[13] [23], \partial_reg[13] [22], 
      \partial_reg[13] [21], \partial_reg[13] [20], \partial_reg[13] [19], 
      \partial_reg[13] [18], \partial_reg[13] [17], \partial_reg[13] [16], 
      \partial_reg[13] [15], \partial_reg[13] [14], \partial_reg[13] [13], 
      \partial_reg[13] [12], \partial_reg[13] [11], \partial_reg[13] [10], 
      \partial_reg[13] [9], \partial_reg[13] [8], \partial_reg[13] [7], 
      \partial_reg[13] [6], \partial_reg[13] [5], \partial_reg[13] [4], 
      \partial_reg[13] [3], \partial_reg[13] [2], \partial_reg[13] [1], 
      \partial_reg[13] [0]}), .s1({uc_32, n_39_350, n_39_349, n_39_348, n_39_347, 
      n_39_346, n_39_345, n_39_344, n_39_343, n_39_342, n_39_341, n_39_340, 
      n_39_339, n_39_338, n_39_337, n_39_336, n_39_335, n_39_334, n_39_333, 
      n_39_332, n_39_331, n_39_330, n_39_329, n_39_328, n_39_327, n_39_326, 
      n_39_325, n_39_324, n_39_323, n_39_322, n_39_321, n_39_320, n_10}), 
      .c1(\c1[11] ));
   PartialAdder__1_1253 genblk1_12_p2 (.a({\partial_reg[13] [31], n_39_350, 
      n_39_349, n_39_348, n_39_347, n_39_346, n_39_345, n_39_344, n_39_343, 
      n_39_342, n_39_341, n_39_340, n_39_339, n_39_338, n_39_337, n_39_336, 
      n_39_335, n_39_334, n_39_333, n_39_332, n_39_331, n_39_330, n_39_329, 
      n_39_328, n_39_327, n_39_326, n_39_325, n_39_324, n_39_323, n_39_322, 
      n_39_321, n_39_320, uc_33}), .b(\c1[11] ), .c({uc_34, 
      \partial_reg[14] [30], \partial_reg[14] [29], \partial_reg[14] [28], 
      \partial_reg[14] [27], \partial_reg[14] [26], \partial_reg[14] [25], 
      \partial_reg[14] [24], \partial_reg[14] [23], \partial_reg[14] [22], 
      \partial_reg[14] [21], \partial_reg[14] [20], \partial_reg[14] [19], 
      \partial_reg[14] [18], \partial_reg[14] [17], \partial_reg[14] [16], 
      \partial_reg[14] [15], \partial_reg[14] [14], \partial_reg[14] [13], 
      \partial_reg[14] [12], \partial_reg[14] [11], \partial_reg[14] [10], 
      \partial_reg[14] [9], \partial_reg[14] [8], \partial_reg[14] [7], 
      \partial_reg[14] [6], \partial_reg[14] [5], \partial_reg[14] [4], 
      \partial_reg[14] [3], \partial_reg[14] [2], \partial_reg[14] [1], 
      \partial_reg[14] [0]}), .s1({uc_35, n_39_382, n_39_381, n_39_380, n_39_379, 
      n_39_378, n_39_377, n_39_376, n_39_375, n_39_374, n_39_373, n_39_372, 
      n_39_371, n_39_370, n_39_369, n_39_368, n_39_367, n_39_366, n_39_365, 
      n_39_364, n_39_363, n_39_362, n_39_361, n_39_360, n_39_359, n_39_358, 
      n_39_357, n_39_356, n_39_355, n_39_354, n_39_353, n_39_352, n_11}), 
      .c1(\c1[12] ));
   PartialAdder__1_1350 genblk1_13_p2 (.a({\partial_reg[14] [31], n_39_382, 
      n_39_381, n_39_380, n_39_379, n_39_378, n_39_377, n_39_376, n_39_375, 
      n_39_374, n_39_373, n_39_372, n_39_371, n_39_370, n_39_369, n_39_368, 
      n_39_367, n_39_366, n_39_365, n_39_364, n_39_363, n_39_362, n_39_361, 
      n_39_360, n_39_359, n_39_358, n_39_357, n_39_356, n_39_355, n_39_354, 
      n_39_353, n_39_352, uc_36}), .b(\c1[12] ), .c({uc_37, 
      \partial_reg[15] [30], \partial_reg[15] [29], \partial_reg[15] [28], 
      \partial_reg[15] [27], \partial_reg[15] [26], \partial_reg[15] [25], 
      \partial_reg[15] [24], \partial_reg[15] [23], \partial_reg[15] [22], 
      \partial_reg[15] [21], \partial_reg[15] [20], \partial_reg[15] [19], 
      \partial_reg[15] [18], \partial_reg[15] [17], \partial_reg[15] [16], 
      \partial_reg[15] [15], \partial_reg[15] [14], \partial_reg[15] [13], 
      \partial_reg[15] [12], \partial_reg[15] [11], \partial_reg[15] [10], 
      \partial_reg[15] [9], \partial_reg[15] [8], \partial_reg[15] [7], 
      \partial_reg[15] [6], \partial_reg[15] [5], \partial_reg[15] [4], 
      \partial_reg[15] [3], \partial_reg[15] [2], \partial_reg[15] [1], 
      \partial_reg[15] [0]}), .s1({uc_38, n_39_414, n_39_413, n_39_412, n_39_411, 
      n_39_410, n_39_409, n_39_408, n_39_407, n_39_406, n_39_405, n_39_404, 
      n_39_403, n_39_402, n_39_401, n_39_400, n_39_399, n_39_398, n_39_397, 
      n_39_396, n_39_395, n_39_394, n_39_393, n_39_392, n_39_391, n_39_390, 
      n_39_389, n_39_388, n_39_387, n_39_386, n_39_385, n_39_384, n_12}), 
      .c1(\c1[13] ));
   PartialAdder__1_1447 genblk1_14_p2 (.a({\partial_reg[15] [31], n_39_414, 
      n_39_413, n_39_412, n_39_411, n_39_410, n_39_409, n_39_408, n_39_407, 
      n_39_406, n_39_405, n_39_404, n_39_403, n_39_402, n_39_401, n_39_400, 
      n_39_399, n_39_398, n_39_397, n_39_396, n_39_395, n_39_394, n_39_393, 
      n_39_392, n_39_391, n_39_390, n_39_389, n_39_388, n_39_387, n_39_386, 
      n_39_385, n_39_384, uc_39}), .b(\c1[13] ), .c({uc_40, 
      \partial_reg[16] [30], \partial_reg[16] [29], \partial_reg[16] [28], 
      \partial_reg[16] [27], \partial_reg[16] [26], \partial_reg[16] [25], 
      \partial_reg[16] [24], \partial_reg[16] [23], \partial_reg[16] [22], 
      \partial_reg[16] [21], \partial_reg[16] [20], \partial_reg[16] [19], 
      \partial_reg[16] [18], \partial_reg[16] [17], \partial_reg[16] [16], 
      \partial_reg[16] [15], \partial_reg[16] [14], \partial_reg[16] [13], 
      \partial_reg[16] [12], \partial_reg[16] [11], \partial_reg[16] [10], 
      \partial_reg[16] [9], \partial_reg[16] [8], \partial_reg[16] [7], 
      \partial_reg[16] [6], \partial_reg[16] [5], \partial_reg[16] [4], 
      \partial_reg[16] [3], \partial_reg[16] [2], \partial_reg[16] [1], 
      \partial_reg[16] [0]}), .s1({uc_41, n_39_446, n_39_445, n_39_444, n_39_443, 
      n_39_442, n_39_441, n_39_440, n_39_439, n_39_438, n_39_437, n_39_436, 
      n_39_435, n_39_434, n_39_433, n_39_432, n_39_431, n_39_430, n_39_429, 
      n_39_428, n_39_427, n_39_426, n_39_425, n_39_424, n_39_423, n_39_422, 
      n_39_421, n_39_420, n_39_419, n_39_418, n_39_417, n_39_416, n_13}), 
      .c1(\c1[14] ));
   PartialAdder__1_1544 genblk1_15_p2 (.a({\partial_reg[16] [31], n_39_446, 
      n_39_445, n_39_444, n_39_443, n_39_442, n_39_441, n_39_440, n_39_439, 
      n_39_438, n_39_437, n_39_436, n_39_435, n_39_434, n_39_433, n_39_432, 
      n_39_431, n_39_430, n_39_429, n_39_428, n_39_427, n_39_426, n_39_425, 
      n_39_424, n_39_423, n_39_422, n_39_421, n_39_420, n_39_419, n_39_418, 
      n_39_417, n_39_416, uc_42}), .b(\c1[14] ), .c({uc_43, 
      \partial_reg[17] [30], \partial_reg[17] [29], \partial_reg[17] [28], 
      \partial_reg[17] [27], \partial_reg[17] [26], \partial_reg[17] [25], 
      \partial_reg[17] [24], \partial_reg[17] [23], \partial_reg[17] [22], 
      \partial_reg[17] [21], \partial_reg[17] [20], \partial_reg[17] [19], 
      \partial_reg[17] [18], \partial_reg[17] [17], \partial_reg[17] [16], 
      \partial_reg[17] [15], \partial_reg[17] [14], \partial_reg[17] [13], 
      \partial_reg[17] [12], \partial_reg[17] [11], \partial_reg[17] [10], 
      \partial_reg[17] [9], \partial_reg[17] [8], \partial_reg[17] [7], 
      \partial_reg[17] [6], \partial_reg[17] [5], \partial_reg[17] [4], 
      \partial_reg[17] [3], \partial_reg[17] [2], \partial_reg[17] [1], 
      \partial_reg[17] [0]}), .s1({uc_44, n_39_478, n_39_477, n_39_476, n_39_475, 
      n_39_474, n_39_473, n_39_472, n_39_471, n_39_470, n_39_469, n_39_468, 
      n_39_467, n_39_466, n_39_465, n_39_464, n_39_463, n_39_462, n_39_461, 
      n_39_460, n_39_459, n_39_458, n_39_457, n_39_456, n_39_455, n_39_454, 
      n_39_453, n_39_452, n_39_451, n_39_450, n_39_449, n_39_448, n_14}), 
      .c1(\c1[15] ));
   PartialAdder__1_1641 genblk1_16_p2 (.a({\partial_reg[17] [31], n_39_478, 
      n_39_477, n_39_476, n_39_475, n_39_474, n_39_473, n_39_472, n_39_471, 
      n_39_470, n_39_469, n_39_468, n_39_467, n_39_466, n_39_465, n_39_464, 
      n_39_463, n_39_462, n_39_461, n_39_460, n_39_459, n_39_458, n_39_457, 
      n_39_456, n_39_455, n_39_454, n_39_453, n_39_452, n_39_451, n_39_450, 
      n_39_449, n_39_448, uc_45}), .b(\c1[15] ), .c({uc_46, 
      \partial_reg[18] [30], \partial_reg[18] [29], \partial_reg[18] [28], 
      \partial_reg[18] [27], \partial_reg[18] [26], \partial_reg[18] [25], 
      \partial_reg[18] [24], \partial_reg[18] [23], \partial_reg[18] [22], 
      \partial_reg[18] [21], \partial_reg[18] [20], \partial_reg[18] [19], 
      \partial_reg[18] [18], \partial_reg[18] [17], \partial_reg[18] [16], 
      \partial_reg[18] [15], \partial_reg[18] [14], \partial_reg[18] [13], 
      \partial_reg[18] [12], \partial_reg[18] [11], \partial_reg[18] [10], 
      \partial_reg[18] [9], \partial_reg[18] [8], \partial_reg[18] [7], 
      \partial_reg[18] [6], \partial_reg[18] [5], \partial_reg[18] [4], 
      \partial_reg[18] [3], \partial_reg[18] [2], \partial_reg[18] [1], 
      \partial_reg[18] [0]}), .s1({uc_47, n_39_510, n_39_509, n_39_508, n_39_507, 
      n_39_506, n_39_505, n_39_504, n_39_503, n_39_502, n_39_501, n_39_500, 
      n_39_499, n_39_498, n_39_497, n_39_496, n_39_495, n_39_494, n_39_493, 
      n_39_492, n_39_491, n_39_490, n_39_489, n_39_488, n_39_487, n_39_486, 
      n_39_485, n_39_484, n_39_483, n_39_482, n_39_481, n_39_480, n_15}), 
      .c1(\c1[16] ));
   PartialAdder__1_1738 genblk1_17_p2 (.a({\partial_reg[18] [31], n_39_510, 
      n_39_509, n_39_508, n_39_507, n_39_506, n_39_505, n_39_504, n_39_503, 
      n_39_502, n_39_501, n_39_500, n_39_499, n_39_498, n_39_497, n_39_496, 
      n_39_495, n_39_494, n_39_493, n_39_492, n_39_491, n_39_490, n_39_489, 
      n_39_488, n_39_487, n_39_486, n_39_485, n_39_484, n_39_483, n_39_482, 
      n_39_481, n_39_480, uc_48}), .b(\c1[16] ), .c({uc_49, 
      \partial_reg[19] [30], \partial_reg[19] [29], \partial_reg[19] [28], 
      \partial_reg[19] [27], \partial_reg[19] [26], \partial_reg[19] [25], 
      \partial_reg[19] [24], \partial_reg[19] [23], \partial_reg[19] [22], 
      \partial_reg[19] [21], \partial_reg[19] [20], \partial_reg[19] [19], 
      \partial_reg[19] [18], \partial_reg[19] [17], \partial_reg[19] [16], 
      \partial_reg[19] [15], \partial_reg[19] [14], \partial_reg[19] [13], 
      \partial_reg[19] [12], \partial_reg[19] [11], \partial_reg[19] [10], 
      \partial_reg[19] [9], \partial_reg[19] [8], \partial_reg[19] [7], 
      \partial_reg[19] [6], \partial_reg[19] [5], \partial_reg[19] [4], 
      \partial_reg[19] [3], \partial_reg[19] [2], \partial_reg[19] [1], 
      \partial_reg[19] [0]}), .s1({uc_50, n_39_542, n_39_541, n_39_540, n_39_539, 
      n_39_538, n_39_537, n_39_536, n_39_535, n_39_534, n_39_533, n_39_532, 
      n_39_531, n_39_530, n_39_529, n_39_528, n_39_527, n_39_526, n_39_525, 
      n_39_524, n_39_523, n_39_522, n_39_521, n_39_520, n_39_519, n_39_518, 
      n_39_517, n_39_516, n_39_515, n_39_514, n_39_513, n_39_512, n_16}), 
      .c1(\c1[17] ));
   PartialAdder__1_1835 genblk1_18_p2 (.a({\partial_reg[19] [31], n_39_542, 
      n_39_541, n_39_540, n_39_539, n_39_538, n_39_537, n_39_536, n_39_535, 
      n_39_534, n_39_533, n_39_532, n_39_531, n_39_530, n_39_529, n_39_528, 
      n_39_527, n_39_526, n_39_525, n_39_524, n_39_523, n_39_522, n_39_521, 
      n_39_520, n_39_519, n_39_518, n_39_517, n_39_516, n_39_515, n_39_514, 
      n_39_513, n_39_512, uc_51}), .b(\c1[17] ), .c({uc_52, 
      \partial_reg[20] [30], \partial_reg[20] [29], \partial_reg[20] [28], 
      \partial_reg[20] [27], \partial_reg[20] [26], \partial_reg[20] [25], 
      \partial_reg[20] [24], \partial_reg[20] [23], \partial_reg[20] [22], 
      \partial_reg[20] [21], \partial_reg[20] [20], \partial_reg[20] [19], 
      \partial_reg[20] [18], \partial_reg[20] [17], \partial_reg[20] [16], 
      \partial_reg[20] [15], \partial_reg[20] [14], \partial_reg[20] [13], 
      \partial_reg[20] [12], \partial_reg[20] [11], \partial_reg[20] [10], 
      \partial_reg[20] [9], \partial_reg[20] [8], \partial_reg[20] [7], 
      \partial_reg[20] [6], \partial_reg[20] [5], \partial_reg[20] [4], 
      \partial_reg[20] [3], \partial_reg[20] [2], \partial_reg[20] [1], 
      \partial_reg[20] [0]}), .s1({uc_53, n_39_574, n_39_573, n_39_572, n_39_571, 
      n_39_570, n_39_569, n_39_568, n_39_567, n_39_566, n_39_565, n_39_564, 
      n_39_563, n_39_562, n_39_561, n_39_560, n_39_559, n_39_558, n_39_557, 
      n_39_556, n_39_555, n_39_554, n_39_553, n_39_552, n_39_551, n_39_550, 
      n_39_549, n_39_548, n_39_547, n_39_546, n_39_545, n_39_544, n_17}), 
      .c1(\c1[18] ));
   PartialAdder__1_1932 genblk1_19_p2 (.a({\partial_reg[20] [31], n_39_574, 
      n_39_573, n_39_572, n_39_571, n_39_570, n_39_569, n_39_568, n_39_567, 
      n_39_566, n_39_565, n_39_564, n_39_563, n_39_562, n_39_561, n_39_560, 
      n_39_559, n_39_558, n_39_557, n_39_556, n_39_555, n_39_554, n_39_553, 
      n_39_552, n_39_551, n_39_550, n_39_549, n_39_548, n_39_547, n_39_546, 
      n_39_545, n_39_544, uc_54}), .b(\c1[18] ), .c({uc_55, 
      \partial_reg[21] [30], \partial_reg[21] [29], \partial_reg[21] [28], 
      \partial_reg[21] [27], \partial_reg[21] [26], \partial_reg[21] [25], 
      \partial_reg[21] [24], \partial_reg[21] [23], \partial_reg[21] [22], 
      \partial_reg[21] [21], \partial_reg[21] [20], \partial_reg[21] [19], 
      \partial_reg[21] [18], \partial_reg[21] [17], \partial_reg[21] [16], 
      \partial_reg[21] [15], \partial_reg[21] [14], \partial_reg[21] [13], 
      \partial_reg[21] [12], \partial_reg[21] [11], \partial_reg[21] [10], 
      \partial_reg[21] [9], \partial_reg[21] [8], \partial_reg[21] [7], 
      \partial_reg[21] [6], \partial_reg[21] [5], \partial_reg[21] [4], 
      \partial_reg[21] [3], \partial_reg[21] [2], \partial_reg[21] [1], 
      \partial_reg[21] [0]}), .s1({uc_56, n_39_606, n_39_605, n_39_604, n_39_603, 
      n_39_602, n_39_601, n_39_600, n_39_599, n_39_598, n_39_597, n_39_596, 
      n_39_595, n_39_594, n_39_593, n_39_592, n_39_591, n_39_590, n_39_589, 
      n_39_588, n_39_587, n_39_586, n_39_585, n_39_584, n_39_583, n_39_582, 
      n_39_581, n_39_580, n_39_579, n_39_578, n_39_577, n_39_576, n_18}), 
      .c1(\c1[19] ));
   PartialAdder__1_2029 genblk1_20_p2 (.a({\partial_reg[21] [31], n_39_606, 
      n_39_605, n_39_604, n_39_603, n_39_602, n_39_601, n_39_600, n_39_599, 
      n_39_598, n_39_597, n_39_596, n_39_595, n_39_594, n_39_593, n_39_592, 
      n_39_591, n_39_590, n_39_589, n_39_588, n_39_587, n_39_586, n_39_585, 
      n_39_584, n_39_583, n_39_582, n_39_581, n_39_580, n_39_579, n_39_578, 
      n_39_577, n_39_576, uc_57}), .b(\c1[19] ), .c({uc_58, 
      \partial_reg[22] [30], \partial_reg[22] [29], \partial_reg[22] [28], 
      \partial_reg[22] [27], \partial_reg[22] [26], \partial_reg[22] [25], 
      \partial_reg[22] [24], \partial_reg[22] [23], \partial_reg[22] [22], 
      \partial_reg[22] [21], \partial_reg[22] [20], \partial_reg[22] [19], 
      \partial_reg[22] [18], \partial_reg[22] [17], \partial_reg[22] [16], 
      \partial_reg[22] [15], \partial_reg[22] [14], \partial_reg[22] [13], 
      \partial_reg[22] [12], \partial_reg[22] [11], \partial_reg[22] [10], 
      \partial_reg[22] [9], \partial_reg[22] [8], \partial_reg[22] [7], 
      \partial_reg[22] [6], \partial_reg[22] [5], \partial_reg[22] [4], 
      \partial_reg[22] [3], \partial_reg[22] [2], \partial_reg[22] [1], 
      \partial_reg[22] [0]}), .s1({uc_59, n_39_638, n_39_637, n_39_636, n_39_635, 
      n_39_634, n_39_633, n_39_632, n_39_631, n_39_630, n_39_629, n_39_628, 
      n_39_627, n_39_626, n_39_625, n_39_624, n_39_623, n_39_622, n_39_621, 
      n_39_620, n_39_619, n_39_618, n_39_617, n_39_616, n_39_615, n_39_614, 
      n_39_613, n_39_612, n_39_611, n_39_610, n_39_609, n_39_608, n_19}), 
      .c1(\c1[20] ));
   PartialAdder__1_2126 genblk1_21_p2 (.a({\partial_reg[22] [31], n_39_638, 
      n_39_637, n_39_636, n_39_635, n_39_634, n_39_633, n_39_632, n_39_631, 
      n_39_630, n_39_629, n_39_628, n_39_627, n_39_626, n_39_625, n_39_624, 
      n_39_623, n_39_622, n_39_621, n_39_620, n_39_619, n_39_618, n_39_617, 
      n_39_616, n_39_615, n_39_614, n_39_613, n_39_612, n_39_611, n_39_610, 
      n_39_609, n_39_608, uc_60}), .b(\c1[20] ), .c({uc_61, 
      \partial_reg[23] [30], \partial_reg[23] [29], \partial_reg[23] [28], 
      \partial_reg[23] [27], \partial_reg[23] [26], \partial_reg[23] [25], 
      \partial_reg[23] [24], \partial_reg[23] [23], \partial_reg[23] [22], 
      \partial_reg[23] [21], \partial_reg[23] [20], \partial_reg[23] [19], 
      \partial_reg[23] [18], \partial_reg[23] [17], \partial_reg[23] [16], 
      \partial_reg[23] [15], \partial_reg[23] [14], \partial_reg[23] [13], 
      \partial_reg[23] [12], \partial_reg[23] [11], \partial_reg[23] [10], 
      \partial_reg[23] [9], \partial_reg[23] [8], \partial_reg[23] [7], 
      \partial_reg[23] [6], \partial_reg[23] [5], \partial_reg[23] [4], 
      \partial_reg[23] [3], \partial_reg[23] [2], \partial_reg[23] [1], 
      \partial_reg[23] [0]}), .s1({uc_62, n_39_670, n_39_669, n_39_668, n_39_667, 
      n_39_666, n_39_665, n_39_664, n_39_663, n_39_662, n_39_661, n_39_660, 
      n_39_659, n_39_658, n_39_657, n_39_656, n_39_655, n_39_654, n_39_653, 
      n_39_652, n_39_651, n_39_650, n_39_649, n_39_648, n_39_647, n_39_646, 
      n_39_645, n_39_644, n_39_643, n_39_642, n_39_641, n_39_640, n_20}), 
      .c1(\c1[21] ));
   PartialAdder__1_2223 genblk1_22_p2 (.a({\partial_reg[23] [31], n_39_670, 
      n_39_669, n_39_668, n_39_667, n_39_666, n_39_665, n_39_664, n_39_663, 
      n_39_662, n_39_661, n_39_660, n_39_659, n_39_658, n_39_657, n_39_656, 
      n_39_655, n_39_654, n_39_653, n_39_652, n_39_651, n_39_650, n_39_649, 
      n_39_648, n_39_647, n_39_646, n_39_645, n_39_644, n_39_643, n_39_642, 
      n_39_641, n_39_640, uc_63}), .b(\c1[21] ), .c({uc_64, 
      \partial_reg[24] [30], \partial_reg[24] [29], \partial_reg[24] [28], 
      \partial_reg[24] [27], \partial_reg[24] [26], \partial_reg[24] [25], 
      \partial_reg[24] [24], \partial_reg[24] [23], \partial_reg[24] [22], 
      \partial_reg[24] [21], \partial_reg[24] [20], \partial_reg[24] [19], 
      \partial_reg[24] [18], \partial_reg[24] [17], \partial_reg[24] [16], 
      \partial_reg[24] [15], \partial_reg[24] [14], \partial_reg[24] [13], 
      \partial_reg[24] [12], \partial_reg[24] [11], \partial_reg[24] [10], 
      \partial_reg[24] [9], \partial_reg[24] [8], \partial_reg[24] [7], 
      \partial_reg[24] [6], \partial_reg[24] [5], \partial_reg[24] [4], 
      \partial_reg[24] [3], \partial_reg[24] [2], \partial_reg[24] [1], 
      \partial_reg[24] [0]}), .s1({uc_65, n_39_702, n_39_701, n_39_700, n_39_699, 
      n_39_698, n_39_697, n_39_696, n_39_695, n_39_694, n_39_693, n_39_692, 
      n_39_691, n_39_690, n_39_689, n_39_688, n_39_687, n_39_686, n_39_685, 
      n_39_684, n_39_683, n_39_682, n_39_681, n_39_680, n_39_679, n_39_678, 
      n_39_677, n_39_676, n_39_675, n_39_674, n_39_673, n_39_672, n_21}), 
      .c1(\c1[22] ));
   PartialAdder__1_2320 genblk1_23_p2 (.a({\partial_reg[24] [31], n_39_702, 
      n_39_701, n_39_700, n_39_699, n_39_698, n_39_697, n_39_696, n_39_695, 
      n_39_694, n_39_693, n_39_692, n_39_691, n_39_690, n_39_689, n_39_688, 
      n_39_687, n_39_686, n_39_685, n_39_684, n_39_683, n_39_682, n_39_681, 
      n_39_680, n_39_679, n_39_678, n_39_677, n_39_676, n_39_675, n_39_674, 
      n_39_673, n_39_672, uc_66}), .b(\c1[22] ), .c({uc_67, 
      \partial_reg[25] [30], \partial_reg[25] [29], \partial_reg[25] [28], 
      \partial_reg[25] [27], \partial_reg[25] [26], \partial_reg[25] [25], 
      \partial_reg[25] [24], \partial_reg[25] [23], \partial_reg[25] [22], 
      \partial_reg[25] [21], \partial_reg[25] [20], \partial_reg[25] [19], 
      \partial_reg[25] [18], \partial_reg[25] [17], \partial_reg[25] [16], 
      \partial_reg[25] [15], \partial_reg[25] [14], \partial_reg[25] [13], 
      \partial_reg[25] [12], \partial_reg[25] [11], \partial_reg[25] [10], 
      \partial_reg[25] [9], \partial_reg[25] [8], \partial_reg[25] [7], 
      \partial_reg[25] [6], \partial_reg[25] [5], \partial_reg[25] [4], 
      \partial_reg[25] [3], \partial_reg[25] [2], \partial_reg[25] [1], 
      \partial_reg[25] [0]}), .s1({uc_68, n_39_734, n_39_733, n_39_732, n_39_731, 
      n_39_730, n_39_729, n_39_728, n_39_727, n_39_726, n_39_725, n_39_724, 
      n_39_723, n_39_722, n_39_721, n_39_720, n_39_719, n_39_718, n_39_717, 
      n_39_716, n_39_715, n_39_714, n_39_713, n_39_712, n_39_711, n_39_710, 
      n_39_709, n_39_708, n_39_707, n_39_706, n_39_705, n_39_704, n_22}), 
      .c1(\c1[23] ));
   PartialAdder__1_2417 genblk1_24_p2 (.a({\partial_reg[25] [31], n_39_734, 
      n_39_733, n_39_732, n_39_731, n_39_730, n_39_729, n_39_728, n_39_727, 
      n_39_726, n_39_725, n_39_724, n_39_723, n_39_722, n_39_721, n_39_720, 
      n_39_719, n_39_718, n_39_717, n_39_716, n_39_715, n_39_714, n_39_713, 
      n_39_712, n_39_711, n_39_710, n_39_709, n_39_708, n_39_707, n_39_706, 
      n_39_705, n_39_704, uc_69}), .b(\c1[23] ), .c({uc_70, 
      \partial_reg[26] [30], \partial_reg[26] [29], \partial_reg[26] [28], 
      \partial_reg[26] [27], \partial_reg[26] [26], \partial_reg[26] [25], 
      \partial_reg[26] [24], \partial_reg[26] [23], \partial_reg[26] [22], 
      \partial_reg[26] [21], \partial_reg[26] [20], \partial_reg[26] [19], 
      \partial_reg[26] [18], \partial_reg[26] [17], \partial_reg[26] [16], 
      \partial_reg[26] [15], \partial_reg[26] [14], \partial_reg[26] [13], 
      \partial_reg[26] [12], \partial_reg[26] [11], \partial_reg[26] [10], 
      \partial_reg[26] [9], \partial_reg[26] [8], \partial_reg[26] [7], 
      \partial_reg[26] [6], \partial_reg[26] [5], \partial_reg[26] [4], 
      \partial_reg[26] [3], \partial_reg[26] [2], \partial_reg[26] [1], 
      \partial_reg[26] [0]}), .s1({uc_71, n_39_766, n_39_765, n_39_764, n_39_763, 
      n_39_762, n_39_761, n_39_760, n_39_759, n_39_758, n_39_757, n_39_756, 
      n_39_755, n_39_754, n_39_753, n_39_752, n_39_751, n_39_750, n_39_749, 
      n_39_748, n_39_747, n_39_746, n_39_745, n_39_744, n_39_743, n_39_742, 
      n_39_741, n_39_740, n_39_739, n_39_738, n_39_737, n_39_736, n_23}), 
      .c1(\c1[24] ));
   PartialAdder__1_2514 genblk1_25_p2 (.a({\partial_reg[26] [31], n_39_766, 
      n_39_765, n_39_764, n_39_763, n_39_762, n_39_761, n_39_760, n_39_759, 
      n_39_758, n_39_757, n_39_756, n_39_755, n_39_754, n_39_753, n_39_752, 
      n_39_751, n_39_750, n_39_749, n_39_748, n_39_747, n_39_746, n_39_745, 
      n_39_744, n_39_743, n_39_742, n_39_741, n_39_740, n_39_739, n_39_738, 
      n_39_737, n_39_736, uc_72}), .b(\c1[24] ), .c({uc_73, 
      \partial_reg[27] [30], \partial_reg[27] [29], \partial_reg[27] [28], 
      \partial_reg[27] [27], \partial_reg[27] [26], \partial_reg[27] [25], 
      \partial_reg[27] [24], \partial_reg[27] [23], \partial_reg[27] [22], 
      \partial_reg[27] [21], \partial_reg[27] [20], \partial_reg[27] [19], 
      \partial_reg[27] [18], \partial_reg[27] [17], \partial_reg[27] [16], 
      \partial_reg[27] [15], \partial_reg[27] [14], \partial_reg[27] [13], 
      \partial_reg[27] [12], \partial_reg[27] [11], \partial_reg[27] [10], 
      \partial_reg[27] [9], \partial_reg[27] [8], \partial_reg[27] [7], 
      \partial_reg[27] [6], \partial_reg[27] [5], \partial_reg[27] [4], 
      \partial_reg[27] [3], \partial_reg[27] [2], \partial_reg[27] [1], 
      \partial_reg[27] [0]}), .s1({uc_74, n_39_798, n_39_797, n_39_796, n_39_795, 
      n_39_794, n_39_793, n_39_792, n_39_791, n_39_790, n_39_789, n_39_788, 
      n_39_787, n_39_786, n_39_785, n_39_784, n_39_783, n_39_782, n_39_781, 
      n_39_780, n_39_779, n_39_778, n_39_777, n_39_776, n_39_775, n_39_774, 
      n_39_773, n_39_772, n_39_771, n_39_770, n_39_769, n_39_768, n_24}), 
      .c1(\c1[25] ));
   PartialAdder__1_2611 genblk1_26_p2 (.a({\partial_reg[27] [31], n_39_798, 
      n_39_797, n_39_796, n_39_795, n_39_794, n_39_793, n_39_792, n_39_791, 
      n_39_790, n_39_789, n_39_788, n_39_787, n_39_786, n_39_785, n_39_784, 
      n_39_783, n_39_782, n_39_781, n_39_780, n_39_779, n_39_778, n_39_777, 
      n_39_776, n_39_775, n_39_774, n_39_773, n_39_772, n_39_771, n_39_770, 
      n_39_769, n_39_768, uc_75}), .b(\c1[25] ), .c({uc_76, 
      \partial_reg[28] [30], \partial_reg[28] [29], \partial_reg[28] [28], 
      \partial_reg[28] [27], \partial_reg[28] [26], \partial_reg[28] [25], 
      \partial_reg[28] [24], \partial_reg[28] [23], \partial_reg[28] [22], 
      \partial_reg[28] [21], \partial_reg[28] [20], \partial_reg[28] [19], 
      \partial_reg[28] [18], \partial_reg[28] [17], \partial_reg[28] [16], 
      \partial_reg[28] [15], \partial_reg[28] [14], \partial_reg[28] [13], 
      \partial_reg[28] [12], \partial_reg[28] [11], \partial_reg[28] [10], 
      \partial_reg[28] [9], \partial_reg[28] [8], \partial_reg[28] [7], 
      \partial_reg[28] [6], \partial_reg[28] [5], \partial_reg[28] [4], 
      \partial_reg[28] [3], \partial_reg[28] [2], \partial_reg[28] [1], 
      \partial_reg[28] [0]}), .s1({uc_77, n_39_830, n_39_829, n_39_828, n_39_827, 
      n_39_826, n_39_825, n_39_824, n_39_823, n_39_822, n_39_821, n_39_820, 
      n_39_819, n_39_818, n_39_817, n_39_816, n_39_815, n_39_814, n_39_813, 
      n_39_812, n_39_811, n_39_810, n_39_809, n_39_808, n_39_807, n_39_806, 
      n_39_805, n_39_804, n_39_803, n_39_802, n_39_801, n_39_800, n_25}), 
      .c1(\c1[26] ));
   PartialAdder__1_2708 genblk1_27_p2 (.a({\partial_reg[28] [31], n_39_830, 
      n_39_829, n_39_828, n_39_827, n_39_826, n_39_825, n_39_824, n_39_823, 
      n_39_822, n_39_821, n_39_820, n_39_819, n_39_818, n_39_817, n_39_816, 
      n_39_815, n_39_814, n_39_813, n_39_812, n_39_811, n_39_810, n_39_809, 
      n_39_808, n_39_807, n_39_806, n_39_805, n_39_804, n_39_803, n_39_802, 
      n_39_801, n_39_800, uc_78}), .b(\c1[26] ), .c({uc_79, 
      \partial_reg[29] [30], \partial_reg[29] [29], \partial_reg[29] [28], 
      \partial_reg[29] [27], \partial_reg[29] [26], \partial_reg[29] [25], 
      \partial_reg[29] [24], \partial_reg[29] [23], \partial_reg[29] [22], 
      \partial_reg[29] [21], \partial_reg[29] [20], \partial_reg[29] [19], 
      \partial_reg[29] [18], \partial_reg[29] [17], \partial_reg[29] [16], 
      \partial_reg[29] [15], \partial_reg[29] [14], \partial_reg[29] [13], 
      \partial_reg[29] [12], \partial_reg[29] [11], \partial_reg[29] [10], 
      \partial_reg[29] [9], \partial_reg[29] [8], \partial_reg[29] [7], 
      \partial_reg[29] [6], \partial_reg[29] [5], \partial_reg[29] [4], 
      \partial_reg[29] [3], \partial_reg[29] [2], \partial_reg[29] [1], 
      \partial_reg[29] [0]}), .s1({uc_80, n_39_862, n_39_861, n_39_860, n_39_859, 
      n_39_858, n_39_857, n_39_856, n_39_855, n_39_854, n_39_853, n_39_852, 
      n_39_851, n_39_850, n_39_849, n_39_848, n_39_847, n_39_846, n_39_845, 
      n_39_844, n_39_843, n_39_842, n_39_841, n_39_840, n_39_839, n_39_838, 
      n_39_837, n_39_836, n_39_835, n_39_834, n_39_833, n_39_832, n_26}), 
      .c1(\c1[27] ));
   PartialAdder__1_2805 genblk1_28_p2 (.a({\partial_reg[29] [31], n_39_862, 
      n_39_861, n_39_860, n_39_859, n_39_858, n_39_857, n_39_856, n_39_855, 
      n_39_854, n_39_853, n_39_852, n_39_851, n_39_850, n_39_849, n_39_848, 
      n_39_847, n_39_846, n_39_845, n_39_844, n_39_843, n_39_842, n_39_841, 
      n_39_840, n_39_839, n_39_838, n_39_837, n_39_836, n_39_835, n_39_834, 
      n_39_833, n_39_832, uc_81}), .b(\c1[27] ), .c({uc_82, 
      \partial_reg[30] [30], \partial_reg[30] [29], \partial_reg[30] [28], 
      \partial_reg[30] [27], \partial_reg[30] [26], \partial_reg[30] [25], 
      \partial_reg[30] [24], \partial_reg[30] [23], \partial_reg[30] [22], 
      \partial_reg[30] [21], \partial_reg[30] [20], \partial_reg[30] [19], 
      \partial_reg[30] [18], \partial_reg[30] [17], \partial_reg[30] [16], 
      \partial_reg[30] [15], \partial_reg[30] [14], \partial_reg[30] [13], 
      \partial_reg[30] [12], \partial_reg[30] [11], \partial_reg[30] [10], 
      \partial_reg[30] [9], \partial_reg[30] [8], \partial_reg[30] [7], 
      \partial_reg[30] [6], \partial_reg[30] [5], \partial_reg[30] [4], 
      \partial_reg[30] [3], \partial_reg[30] [2], \partial_reg[30] [1], 
      \partial_reg[30] [0]}), .s1({uc_83, n_39_863, n_39_831, n_39_799, n_39_767, 
      n_39_735, n_39_703, n_39_671, n_39_639, n_39_607, n_39_575, n_39_543, 
      n_39_511, n_39_479, n_39_447, n_39_415, n_39_383, n_39_351, n_39_319, 
      n_39_287, n_39_255, n_39_223, n_39_191, n_39_159, n_39_127, n_39_95, 
      n_39_63, n_39_31, n_39_867, n_39_866, n_39_865, n_39_864, n_27}), .c1(
      \c1[28] ));
   PartialAdder__0_47 genblk1_29_p2 (.a({\partial_reg[30] [31], n_39_863, 
      n_39_831, n_39_799, n_39_767, n_39_735, n_39_703, n_39_671, n_39_639, 
      n_39_607, n_39_575, n_39_543, n_39_511, n_39_479, n_39_447, n_39_415, 
      n_39_383, n_39_351, n_39_319, n_39_287, n_39_255, n_39_223, n_39_191, 
      n_39_159, n_39_127, n_39_95, n_39_63, n_39_31, n_39_867, n_39_866, 
      n_39_865, n_39_864, uc_84}), .b(\c1[28] ), .c({uc_85, 
      \partial_reg[31] [30], \partial_reg[31] [29], \partial_reg[31] [28], 
      \partial_reg[31] [27], \partial_reg[31] [26], \partial_reg[31] [25], 
      \partial_reg[31] [24], \partial_reg[31] [23], \partial_reg[31] [22], 
      \partial_reg[31] [21], \partial_reg[31] [20], \partial_reg[31] [19], 
      \partial_reg[31] [18], \partial_reg[31] [17], \partial_reg[31] [16], 
      \partial_reg[31] [15], \partial_reg[31] [14], \partial_reg[31] [13], 
      \partial_reg[31] [12], \partial_reg[31] [11], \partial_reg[31] [10], 
      \partial_reg[31] [9], \partial_reg[31] [8], \partial_reg[31] [7], 
      \partial_reg[31] [6], \partial_reg[31] [5], \partial_reg[31] [4], 
      \partial_reg[31] [3], \partial_reg[31] [2], \partial_reg[31] [1], 
      \partial_reg[31] [0]}), .s1({uc_86, \s1[29] [31], \s1[29] [30], 
      \s1[29] [29], \s1[29] [28], \s1[29] [27], \s1[29] [26], \s1[29] [25], 
      \s1[29] [24], \s1[29] [23], \s1[29] [22], \s1[29] [21], \s1[29] [20], 
      \s1[29] [19], \s1[29] [18], \s1[29] [17], \s1[29] [16], \s1[29] [15], 
      \s1[29] [14], \s1[29] [13], \s1[29] [12], \s1[29] [11], \s1[29] [10], 
      \s1[29] [9], \s1[29] [8], \s1[29] [7], \s1[29] [6], \s1[29] [5], 
      \s1[29] [4], \s1[29] [3], \s1[29] [2], \s1[29] [1], \s1[29] [0]}), 
      .c1(\c1[29] ));
   adderPlus final (.a({\partial_reg[31] [31], \s1[29] [31], \s1[29] [30], 
      \s1[29] [29], \s1[29] [28], \s1[29] [27], \s1[29] [26], \s1[29] [25], 
      \s1[29] [24], \s1[29] [23], \s1[29] [22], \s1[29] [21], \s1[29] [20], 
      \s1[29] [19], \s1[29] [18], \s1[29] [17], \s1[29] [16], \s1[29] [15], 
      \s1[29] [14], \s1[29] [13], \s1[29] [12], \s1[29] [11], \s1[29] [10], 
      \s1[29] [9], \s1[29] [8], \s1[29] [7], \s1[29] [6], \s1[29] [5], 
      \s1[29] [4], \s1[29] [3], \s1[29] [2], \s1[29] [1]}), .b(\c1[29] ), 
      .sum({n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
      n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, 
      n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29}), .cout(n_28));
   INV_X1 i_4_0_1 (.A(a[0]), .ZN(n_4_0_1));
   NOR2_X1 i_4_0_2 (.A1(n_4_0_0), .A2(n_4_0_1), .ZN(out[0]));
   INV_X1 i_4_0_3 (.A(op1[1]), .ZN(n_4_0_2));
   NOR2_X1 i_4_0_4 (.A1(n_4_0_0), .A2(n_4_0_2), .ZN(\partial_reg[0] [1]));
   INV_X1 i_4_0_5 (.A(op1[2]), .ZN(n_4_0_3));
   NOR2_X1 i_4_0_6 (.A1(n_4_0_0), .A2(n_4_0_3), .ZN(\partial_reg[0] [2]));
   INV_X1 i_4_0_7 (.A(op1[3]), .ZN(n_4_0_4));
   NOR2_X1 i_4_0_8 (.A1(n_4_0_0), .A2(n_4_0_4), .ZN(\partial_reg[0] [3]));
   INV_X1 i_4_0_9 (.A(op1[4]), .ZN(n_4_0_5));
   NOR2_X1 i_4_0_10 (.A1(n_4_0_0), .A2(n_4_0_5), .ZN(\partial_reg[0] [4]));
   INV_X1 i_4_0_11 (.A(op1[5]), .ZN(n_4_0_6));
   NOR2_X1 i_4_0_12 (.A1(n_4_0_0), .A2(n_4_0_6), .ZN(\partial_reg[0] [5]));
   INV_X1 i_4_0_13 (.A(op1[6]), .ZN(n_4_0_7));
   NOR2_X1 i_4_0_14 (.A1(n_4_0_0), .A2(n_4_0_7), .ZN(\partial_reg[0] [6]));
   INV_X1 i_4_0_15 (.A(op1[7]), .ZN(n_4_0_8));
   NOR2_X1 i_4_0_16 (.A1(n_4_0_0), .A2(n_4_0_8), .ZN(\partial_reg[0] [7]));
   INV_X1 i_4_0_17 (.A(op1[8]), .ZN(n_4_0_9));
   NOR2_X1 i_4_0_18 (.A1(n_4_0_0), .A2(n_4_0_9), .ZN(\partial_reg[0] [8]));
   INV_X1 i_4_0_19 (.A(op1[9]), .ZN(n_4_0_10));
   NOR2_X1 i_4_0_20 (.A1(n_4_0_0), .A2(n_4_0_10), .ZN(\partial_reg[0] [9]));
   INV_X1 i_4_0_21 (.A(op1[10]), .ZN(n_4_0_11));
   NOR2_X1 i_4_0_22 (.A1(n_4_0_0), .A2(n_4_0_11), .ZN(\partial_reg[0] [10]));
   INV_X1 i_4_0_23 (.A(op1[11]), .ZN(n_4_0_12));
   NOR2_X1 i_4_0_24 (.A1(n_4_0_0), .A2(n_4_0_12), .ZN(\partial_reg[0] [11]));
   INV_X1 i_4_0_25 (.A(op1[12]), .ZN(n_4_0_13));
   NOR2_X1 i_4_0_26 (.A1(n_4_0_0), .A2(n_4_0_13), .ZN(\partial_reg[0] [12]));
   INV_X1 i_4_0_27 (.A(op1[13]), .ZN(n_4_0_14));
   NOR2_X1 i_4_0_28 (.A1(n_4_0_0), .A2(n_4_0_14), .ZN(\partial_reg[0] [13]));
   INV_X1 i_4_0_29 (.A(op1[14]), .ZN(n_4_0_15));
   NOR2_X1 i_4_0_30 (.A1(n_4_0_0), .A2(n_4_0_15), .ZN(\partial_reg[0] [14]));
   INV_X1 i_4_0_31 (.A(op1[15]), .ZN(n_4_0_16));
   NOR2_X1 i_4_0_32 (.A1(n_4_0_0), .A2(n_4_0_16), .ZN(\partial_reg[0] [15]));
   INV_X1 i_4_0_33 (.A(op1[16]), .ZN(n_4_0_17));
   NOR2_X1 i_4_0_34 (.A1(n_4_0_0), .A2(n_4_0_17), .ZN(\partial_reg[0] [16]));
   INV_X1 i_4_0_35 (.A(op1[17]), .ZN(n_4_0_18));
   NOR2_X1 i_4_0_36 (.A1(n_4_0_0), .A2(n_4_0_18), .ZN(\partial_reg[0] [17]));
   INV_X1 i_4_0_37 (.A(op1[18]), .ZN(n_4_0_19));
   NOR2_X1 i_4_0_38 (.A1(n_4_0_0), .A2(n_4_0_19), .ZN(\partial_reg[0] [18]));
   INV_X1 i_4_0_39 (.A(op1[19]), .ZN(n_4_0_20));
   NOR2_X1 i_4_0_40 (.A1(n_4_0_0), .A2(n_4_0_20), .ZN(\partial_reg[0] [19]));
   INV_X1 i_4_0_41 (.A(op1[20]), .ZN(n_4_0_21));
   NOR2_X1 i_4_0_42 (.A1(n_4_0_0), .A2(n_4_0_21), .ZN(\partial_reg[0] [20]));
   INV_X1 i_4_0_43 (.A(op1[21]), .ZN(n_4_0_22));
   NOR2_X1 i_4_0_44 (.A1(n_4_0_0), .A2(n_4_0_22), .ZN(\partial_reg[0] [21]));
   INV_X1 i_4_0_45 (.A(op1[22]), .ZN(n_4_0_23));
   NOR2_X1 i_4_0_46 (.A1(n_4_0_0), .A2(n_4_0_23), .ZN(\partial_reg[0] [22]));
   INV_X1 i_4_0_47 (.A(op1[23]), .ZN(n_4_0_24));
   NOR2_X1 i_4_0_48 (.A1(n_4_0_0), .A2(n_4_0_24), .ZN(\partial_reg[0] [23]));
   INV_X1 i_4_0_49 (.A(op1[24]), .ZN(n_4_0_25));
   NOR2_X1 i_4_0_50 (.A1(n_4_0_0), .A2(n_4_0_25), .ZN(\partial_reg[0] [24]));
   INV_X1 i_4_0_51 (.A(op1[25]), .ZN(n_4_0_26));
   NOR2_X1 i_4_0_52 (.A1(n_4_0_0), .A2(n_4_0_26), .ZN(\partial_reg[0] [25]));
   INV_X1 i_4_0_53 (.A(op1[26]), .ZN(n_4_0_27));
   NOR2_X1 i_4_0_54 (.A1(n_4_0_0), .A2(n_4_0_27), .ZN(\partial_reg[0] [26]));
   INV_X1 i_4_0_55 (.A(op1[27]), .ZN(n_4_0_28));
   NOR2_X1 i_4_0_56 (.A1(n_4_0_0), .A2(n_4_0_28), .ZN(\partial_reg[0] [27]));
   INV_X1 i_4_0_57 (.A(op1[28]), .ZN(n_4_0_29));
   NOR2_X1 i_4_0_58 (.A1(n_4_0_0), .A2(n_4_0_29), .ZN(\partial_reg[0] [28]));
   NOR2_X1 i_4_0_60 (.A1(n_4_0_0), .A2(n_4_0_30), .ZN(\partial_reg[0] [29]));
   NOR2_X1 i_4_0_62 (.A1(n_4_0_0), .A2(n_4_0_31), .ZN(\partial_reg[0] [30]));
   NOR2_X1 i_4_0_66 (.A1(n_4_0_33), .A2(n_4_0_1), .ZN(\partial_reg[1] [0]));
   NOR2_X1 i_4_0_67 (.A1(n_4_0_33), .A2(n_4_0_2), .ZN(\partial_reg[1] [1]));
   NOR2_X1 i_4_0_68 (.A1(n_4_0_33), .A2(n_4_0_3), .ZN(\partial_reg[1] [2]));
   NOR2_X1 i_4_0_69 (.A1(n_4_0_33), .A2(n_4_0_4), .ZN(\partial_reg[1] [3]));
   NOR2_X1 i_4_0_70 (.A1(n_4_0_33), .A2(n_4_0_5), .ZN(\partial_reg[1] [4]));
   NOR2_X1 i_4_0_71 (.A1(n_4_0_33), .A2(n_4_0_6), .ZN(\partial_reg[1] [5]));
   NOR2_X1 i_4_0_72 (.A1(n_4_0_33), .A2(n_4_0_7), .ZN(\partial_reg[1] [6]));
   NOR2_X1 i_4_0_73 (.A1(n_4_0_33), .A2(n_4_0_8), .ZN(\partial_reg[1] [7]));
   NOR2_X1 i_4_0_74 (.A1(n_4_0_33), .A2(n_4_0_9), .ZN(\partial_reg[1] [8]));
   NOR2_X1 i_4_0_75 (.A1(n_4_0_33), .A2(n_4_0_10), .ZN(\partial_reg[1] [9]));
   NOR2_X1 i_4_0_76 (.A1(n_4_0_33), .A2(n_4_0_11), .ZN(\partial_reg[1] [10]));
   NOR2_X1 i_4_0_77 (.A1(n_4_0_33), .A2(n_4_0_12), .ZN(\partial_reg[1] [11]));
   NOR2_X1 i_4_0_78 (.A1(n_4_0_33), .A2(n_4_0_13), .ZN(\partial_reg[1] [12]));
   NOR2_X1 i_4_0_79 (.A1(n_4_0_33), .A2(n_4_0_14), .ZN(\partial_reg[1] [13]));
   NOR2_X1 i_4_0_80 (.A1(n_4_0_33), .A2(n_4_0_15), .ZN(\partial_reg[1] [14]));
   NOR2_X1 i_4_0_81 (.A1(n_4_0_33), .A2(n_4_0_16), .ZN(\partial_reg[1] [15]));
   NOR2_X1 i_4_0_82 (.A1(n_4_0_33), .A2(n_4_0_17), .ZN(\partial_reg[1] [16]));
   NOR2_X1 i_4_0_83 (.A1(n_4_0_33), .A2(n_4_0_18), .ZN(\partial_reg[1] [17]));
   NOR2_X1 i_4_0_84 (.A1(n_4_0_33), .A2(n_4_0_19), .ZN(\partial_reg[1] [18]));
   NOR2_X1 i_4_0_85 (.A1(n_4_0_33), .A2(n_4_0_20), .ZN(\partial_reg[1] [19]));
   NOR2_X1 i_4_0_86 (.A1(n_4_0_33), .A2(n_4_0_21), .ZN(\partial_reg[1] [20]));
   NOR2_X1 i_4_0_87 (.A1(n_4_0_33), .A2(n_4_0_22), .ZN(\partial_reg[1] [21]));
   NOR2_X1 i_4_0_88 (.A1(n_4_0_33), .A2(n_4_0_23), .ZN(\partial_reg[1] [22]));
   NOR2_X1 i_4_0_89 (.A1(n_4_0_33), .A2(n_4_0_24), .ZN(\partial_reg[1] [23]));
   NOR2_X1 i_4_0_90 (.A1(n_4_0_33), .A2(n_4_0_25), .ZN(\partial_reg[1] [24]));
   NOR2_X1 i_4_0_91 (.A1(n_4_0_33), .A2(n_4_0_26), .ZN(\partial_reg[1] [25]));
   NOR2_X1 i_4_0_92 (.A1(n_4_0_33), .A2(n_4_0_27), .ZN(\partial_reg[1] [26]));
   NOR2_X1 i_4_0_93 (.A1(n_4_0_33), .A2(n_4_0_28), .ZN(\partial_reg[1] [27]));
   NOR2_X1 i_4_0_94 (.A1(n_4_0_33), .A2(n_4_0_29), .ZN(\partial_reg[1] [28]));
   NOR2_X1 i_4_0_95 (.A1(n_4_0_33), .A2(n_4_0_30), .ZN(\partial_reg[1] [29]));
   NOR2_X1 i_4_0_99 (.A1(n_4_0_34), .A2(n_4_0_1), .ZN(\partial_reg[2] [0]));
   NOR2_X1 i_4_0_100 (.A1(n_4_0_34), .A2(n_4_0_2), .ZN(\partial_reg[2] [1]));
   NOR2_X1 i_4_0_101 (.A1(n_4_0_34), .A2(n_4_0_3), .ZN(\partial_reg[2] [2]));
   NOR2_X1 i_4_0_102 (.A1(n_4_0_34), .A2(n_4_0_4), .ZN(\partial_reg[2] [3]));
   NOR2_X1 i_4_0_103 (.A1(n_4_0_34), .A2(n_4_0_5), .ZN(\partial_reg[2] [4]));
   NOR2_X1 i_4_0_104 (.A1(n_4_0_34), .A2(n_4_0_6), .ZN(\partial_reg[2] [5]));
   NOR2_X1 i_4_0_105 (.A1(n_4_0_34), .A2(n_4_0_7), .ZN(\partial_reg[2] [6]));
   NOR2_X1 i_4_0_106 (.A1(n_4_0_34), .A2(n_4_0_8), .ZN(\partial_reg[2] [7]));
   NOR2_X1 i_4_0_107 (.A1(n_4_0_34), .A2(n_4_0_9), .ZN(\partial_reg[2] [8]));
   NOR2_X1 i_4_0_108 (.A1(n_4_0_34), .A2(n_4_0_10), .ZN(\partial_reg[2] [9]));
   NOR2_X1 i_4_0_109 (.A1(n_4_0_34), .A2(n_4_0_11), .ZN(\partial_reg[2] [10]));
   NOR2_X1 i_4_0_110 (.A1(n_4_0_34), .A2(n_4_0_12), .ZN(\partial_reg[2] [11]));
   NOR2_X1 i_4_0_111 (.A1(n_4_0_34), .A2(n_4_0_13), .ZN(\partial_reg[2] [12]));
   NOR2_X1 i_4_0_112 (.A1(n_4_0_34), .A2(n_4_0_14), .ZN(\partial_reg[2] [13]));
   NOR2_X1 i_4_0_113 (.A1(n_4_0_34), .A2(n_4_0_15), .ZN(\partial_reg[2] [14]));
   NOR2_X1 i_4_0_114 (.A1(n_4_0_34), .A2(n_4_0_16), .ZN(\partial_reg[2] [15]));
   NOR2_X1 i_4_0_115 (.A1(n_4_0_34), .A2(n_4_0_17), .ZN(\partial_reg[2] [16]));
   NOR2_X1 i_4_0_116 (.A1(n_4_0_34), .A2(n_4_0_18), .ZN(\partial_reg[2] [17]));
   NOR2_X1 i_4_0_117 (.A1(n_4_0_34), .A2(n_4_0_19), .ZN(\partial_reg[2] [18]));
   NOR2_X1 i_4_0_118 (.A1(n_4_0_34), .A2(n_4_0_20), .ZN(\partial_reg[2] [19]));
   NOR2_X1 i_4_0_119 (.A1(n_4_0_34), .A2(n_4_0_21), .ZN(\partial_reg[2] [20]));
   NOR2_X1 i_4_0_120 (.A1(n_4_0_34), .A2(n_4_0_22), .ZN(\partial_reg[2] [21]));
   NOR2_X1 i_4_0_121 (.A1(n_4_0_34), .A2(n_4_0_23), .ZN(\partial_reg[2] [22]));
   NOR2_X1 i_4_0_122 (.A1(n_4_0_34), .A2(n_4_0_24), .ZN(\partial_reg[2] [23]));
   NOR2_X1 i_4_0_123 (.A1(n_4_0_34), .A2(n_4_0_25), .ZN(\partial_reg[2] [24]));
   NOR2_X1 i_4_0_124 (.A1(n_4_0_34), .A2(n_4_0_26), .ZN(\partial_reg[2] [25]));
   NOR2_X1 i_4_0_125 (.A1(n_4_0_34), .A2(n_4_0_27), .ZN(\partial_reg[2] [26]));
   NOR2_X1 i_4_0_126 (.A1(n_4_0_34), .A2(n_4_0_28), .ZN(\partial_reg[2] [27]));
   NOR2_X1 i_4_0_127 (.A1(n_4_0_34), .A2(n_4_0_29), .ZN(\partial_reg[2] [28]));
   NOR2_X1 i_4_0_130 (.A1(n_4_0_34), .A2(n_4_0_32), .ZN(\partial_reg[2] [31]));
   INV_X1 i_4_0_131 (.A(op2[3]), .ZN(n_4_0_35));
   NOR2_X1 i_4_0_132 (.A1(n_4_0_35), .A2(n_4_0_1), .ZN(\partial_reg[3] [0]));
   NOR2_X1 i_4_0_133 (.A1(n_4_0_35), .A2(n_4_0_2), .ZN(\partial_reg[3] [1]));
   NOR2_X1 i_4_0_134 (.A1(n_4_0_35), .A2(n_4_0_3), .ZN(\partial_reg[3] [2]));
   NOR2_X1 i_4_0_135 (.A1(n_4_0_35), .A2(n_4_0_4), .ZN(\partial_reg[3] [3]));
   NOR2_X1 i_4_0_136 (.A1(n_4_0_35), .A2(n_4_0_5), .ZN(\partial_reg[3] [4]));
   NOR2_X1 i_4_0_137 (.A1(n_4_0_35), .A2(n_4_0_6), .ZN(\partial_reg[3] [5]));
   NOR2_X1 i_4_0_138 (.A1(n_4_0_35), .A2(n_4_0_7), .ZN(\partial_reg[3] [6]));
   NOR2_X1 i_4_0_139 (.A1(n_4_0_35), .A2(n_4_0_8), .ZN(\partial_reg[3] [7]));
   NOR2_X1 i_4_0_140 (.A1(n_4_0_35), .A2(n_4_0_9), .ZN(\partial_reg[3] [8]));
   NOR2_X1 i_4_0_141 (.A1(n_4_0_35), .A2(n_4_0_10), .ZN(\partial_reg[3] [9]));
   NOR2_X1 i_4_0_142 (.A1(n_4_0_35), .A2(n_4_0_11), .ZN(\partial_reg[3] [10]));
   NOR2_X1 i_4_0_143 (.A1(n_4_0_35), .A2(n_4_0_12), .ZN(\partial_reg[3] [11]));
   NOR2_X1 i_4_0_144 (.A1(n_4_0_35), .A2(n_4_0_13), .ZN(\partial_reg[3] [12]));
   NOR2_X1 i_4_0_145 (.A1(n_4_0_35), .A2(n_4_0_14), .ZN(\partial_reg[3] [13]));
   NOR2_X1 i_4_0_146 (.A1(n_4_0_35), .A2(n_4_0_15), .ZN(\partial_reg[3] [14]));
   NOR2_X1 i_4_0_147 (.A1(n_4_0_35), .A2(n_4_0_16), .ZN(\partial_reg[3] [15]));
   NOR2_X1 i_4_0_148 (.A1(n_4_0_35), .A2(n_4_0_17), .ZN(\partial_reg[3] [16]));
   NOR2_X1 i_4_0_149 (.A1(n_4_0_35), .A2(n_4_0_18), .ZN(\partial_reg[3] [17]));
   NOR2_X1 i_4_0_150 (.A1(n_4_0_35), .A2(n_4_0_19), .ZN(\partial_reg[3] [18]));
   NOR2_X1 i_4_0_151 (.A1(n_4_0_35), .A2(n_4_0_20), .ZN(\partial_reg[3] [19]));
   NOR2_X1 i_4_0_152 (.A1(n_4_0_35), .A2(n_4_0_21), .ZN(\partial_reg[3] [20]));
   NOR2_X1 i_4_0_153 (.A1(n_4_0_35), .A2(n_4_0_22), .ZN(\partial_reg[3] [21]));
   NOR2_X1 i_4_0_154 (.A1(n_4_0_35), .A2(n_4_0_23), .ZN(\partial_reg[3] [22]));
   NOR2_X1 i_4_0_155 (.A1(n_4_0_35), .A2(n_4_0_24), .ZN(\partial_reg[3] [23]));
   NOR2_X1 i_4_0_156 (.A1(n_4_0_35), .A2(n_4_0_25), .ZN(\partial_reg[3] [24]));
   NOR2_X1 i_4_0_157 (.A1(n_4_0_35), .A2(n_4_0_26), .ZN(\partial_reg[3] [25]));
   NOR2_X1 i_4_0_158 (.A1(n_4_0_35), .A2(n_4_0_27), .ZN(\partial_reg[3] [26]));
   NOR2_X1 i_4_0_159 (.A1(n_4_0_35), .A2(n_4_0_28), .ZN(\partial_reg[3] [27]));
   NOR2_X1 i_4_0_160 (.A1(n_4_0_35), .A2(n_4_0_29), .ZN(\partial_reg[3] [28]));
   NOR2_X1 i_4_0_161 (.A1(n_4_0_35), .A2(n_4_0_30), .ZN(\partial_reg[3] [29]));
   NOR2_X1 i_4_0_162 (.A1(n_4_0_35), .A2(n_4_0_31), .ZN(\partial_reg[3] [30]));
   NOR2_X1 i_4_0_163 (.A1(n_4_0_35), .A2(n_4_0_32), .ZN(\partial_reg[3] [31]));
   INV_X1 i_4_0_164 (.A(op2[4]), .ZN(n_4_0_36));
   NOR2_X1 i_4_0_165 (.A1(n_4_0_36), .A2(n_4_0_1), .ZN(\partial_reg[4] [0]));
   NOR2_X1 i_4_0_166 (.A1(n_4_0_36), .A2(n_4_0_2), .ZN(\partial_reg[4] [1]));
   NOR2_X1 i_4_0_167 (.A1(n_4_0_36), .A2(n_4_0_3), .ZN(\partial_reg[4] [2]));
   NOR2_X1 i_4_0_168 (.A1(n_4_0_36), .A2(n_4_0_4), .ZN(\partial_reg[4] [3]));
   NOR2_X1 i_4_0_169 (.A1(n_4_0_36), .A2(n_4_0_5), .ZN(\partial_reg[4] [4]));
   NOR2_X1 i_4_0_170 (.A1(n_4_0_36), .A2(n_4_0_6), .ZN(\partial_reg[4] [5]));
   NOR2_X1 i_4_0_171 (.A1(n_4_0_36), .A2(n_4_0_7), .ZN(\partial_reg[4] [6]));
   NOR2_X1 i_4_0_172 (.A1(n_4_0_36), .A2(n_4_0_8), .ZN(\partial_reg[4] [7]));
   NOR2_X1 i_4_0_173 (.A1(n_4_0_36), .A2(n_4_0_9), .ZN(\partial_reg[4] [8]));
   NOR2_X1 i_4_0_174 (.A1(n_4_0_36), .A2(n_4_0_10), .ZN(\partial_reg[4] [9]));
   NOR2_X1 i_4_0_175 (.A1(n_4_0_36), .A2(n_4_0_11), .ZN(\partial_reg[4] [10]));
   NOR2_X1 i_4_0_176 (.A1(n_4_0_36), .A2(n_4_0_12), .ZN(\partial_reg[4] [11]));
   NOR2_X1 i_4_0_177 (.A1(n_4_0_36), .A2(n_4_0_13), .ZN(\partial_reg[4] [12]));
   NOR2_X1 i_4_0_178 (.A1(n_4_0_36), .A2(n_4_0_14), .ZN(\partial_reg[4] [13]));
   NOR2_X1 i_4_0_179 (.A1(n_4_0_36), .A2(n_4_0_15), .ZN(\partial_reg[4] [14]));
   NOR2_X1 i_4_0_180 (.A1(n_4_0_36), .A2(n_4_0_16), .ZN(\partial_reg[4] [15]));
   NOR2_X1 i_4_0_181 (.A1(n_4_0_36), .A2(n_4_0_17), .ZN(\partial_reg[4] [16]));
   NOR2_X1 i_4_0_182 (.A1(n_4_0_36), .A2(n_4_0_18), .ZN(\partial_reg[4] [17]));
   NOR2_X1 i_4_0_183 (.A1(n_4_0_36), .A2(n_4_0_19), .ZN(\partial_reg[4] [18]));
   NOR2_X1 i_4_0_184 (.A1(n_4_0_36), .A2(n_4_0_20), .ZN(\partial_reg[4] [19]));
   NOR2_X1 i_4_0_185 (.A1(n_4_0_36), .A2(n_4_0_21), .ZN(\partial_reg[4] [20]));
   NOR2_X1 i_4_0_186 (.A1(n_4_0_36), .A2(n_4_0_22), .ZN(\partial_reg[4] [21]));
   NOR2_X1 i_4_0_187 (.A1(n_4_0_36), .A2(n_4_0_23), .ZN(\partial_reg[4] [22]));
   NOR2_X1 i_4_0_188 (.A1(n_4_0_36), .A2(n_4_0_24), .ZN(\partial_reg[4] [23]));
   NOR2_X1 i_4_0_189 (.A1(n_4_0_36), .A2(n_4_0_25), .ZN(\partial_reg[4] [24]));
   NOR2_X1 i_4_0_190 (.A1(n_4_0_36), .A2(n_4_0_26), .ZN(\partial_reg[4] [25]));
   NOR2_X1 i_4_0_191 (.A1(n_4_0_36), .A2(n_4_0_27), .ZN(\partial_reg[4] [26]));
   NOR2_X1 i_4_0_192 (.A1(n_4_0_36), .A2(n_4_0_28), .ZN(\partial_reg[4] [27]));
   NOR2_X1 i_4_0_193 (.A1(n_4_0_36), .A2(n_4_0_29), .ZN(\partial_reg[4] [28]));
   NOR2_X1 i_4_0_194 (.A1(n_4_0_36), .A2(n_4_0_30), .ZN(\partial_reg[4] [29]));
   NOR2_X1 i_4_0_195 (.A1(n_4_0_36), .A2(n_4_0_31), .ZN(\partial_reg[4] [30]));
   NOR2_X1 i_4_0_196 (.A1(n_4_0_36), .A2(n_4_0_32), .ZN(\partial_reg[4] [31]));
   INV_X1 i_4_0_197 (.A(op2[5]), .ZN(n_4_0_37));
   NOR2_X1 i_4_0_198 (.A1(n_4_0_37), .A2(n_4_0_1), .ZN(\partial_reg[5] [0]));
   NOR2_X1 i_4_0_199 (.A1(n_4_0_37), .A2(n_4_0_2), .ZN(\partial_reg[5] [1]));
   NOR2_X1 i_4_0_200 (.A1(n_4_0_37), .A2(n_4_0_3), .ZN(\partial_reg[5] [2]));
   NOR2_X1 i_4_0_201 (.A1(n_4_0_37), .A2(n_4_0_4), .ZN(\partial_reg[5] [3]));
   NOR2_X1 i_4_0_202 (.A1(n_4_0_37), .A2(n_4_0_5), .ZN(\partial_reg[5] [4]));
   NOR2_X1 i_4_0_203 (.A1(n_4_0_37), .A2(n_4_0_6), .ZN(\partial_reg[5] [5]));
   NOR2_X1 i_4_0_204 (.A1(n_4_0_37), .A2(n_4_0_7), .ZN(\partial_reg[5] [6]));
   NOR2_X1 i_4_0_205 (.A1(n_4_0_37), .A2(n_4_0_8), .ZN(\partial_reg[5] [7]));
   NOR2_X1 i_4_0_206 (.A1(n_4_0_37), .A2(n_4_0_9), .ZN(\partial_reg[5] [8]));
   NOR2_X1 i_4_0_207 (.A1(n_4_0_37), .A2(n_4_0_10), .ZN(\partial_reg[5] [9]));
   NOR2_X1 i_4_0_208 (.A1(n_4_0_37), .A2(n_4_0_11), .ZN(\partial_reg[5] [10]));
   NOR2_X1 i_4_0_209 (.A1(n_4_0_37), .A2(n_4_0_12), .ZN(\partial_reg[5] [11]));
   NOR2_X1 i_4_0_210 (.A1(n_4_0_37), .A2(n_4_0_13), .ZN(\partial_reg[5] [12]));
   NOR2_X1 i_4_0_211 (.A1(n_4_0_37), .A2(n_4_0_14), .ZN(\partial_reg[5] [13]));
   NOR2_X1 i_4_0_212 (.A1(n_4_0_37), .A2(n_4_0_15), .ZN(\partial_reg[5] [14]));
   NOR2_X1 i_4_0_213 (.A1(n_4_0_37), .A2(n_4_0_16), .ZN(\partial_reg[5] [15]));
   NOR2_X1 i_4_0_214 (.A1(n_4_0_37), .A2(n_4_0_17), .ZN(\partial_reg[5] [16]));
   NOR2_X1 i_4_0_215 (.A1(n_4_0_37), .A2(n_4_0_18), .ZN(\partial_reg[5] [17]));
   NOR2_X1 i_4_0_216 (.A1(n_4_0_37), .A2(n_4_0_19), .ZN(\partial_reg[5] [18]));
   NOR2_X1 i_4_0_217 (.A1(n_4_0_37), .A2(n_4_0_20), .ZN(\partial_reg[5] [19]));
   NOR2_X1 i_4_0_218 (.A1(n_4_0_37), .A2(n_4_0_21), .ZN(\partial_reg[5] [20]));
   NOR2_X1 i_4_0_219 (.A1(n_4_0_37), .A2(n_4_0_22), .ZN(\partial_reg[5] [21]));
   NOR2_X1 i_4_0_220 (.A1(n_4_0_37), .A2(n_4_0_23), .ZN(\partial_reg[5] [22]));
   NOR2_X1 i_4_0_221 (.A1(n_4_0_37), .A2(n_4_0_24), .ZN(\partial_reg[5] [23]));
   NOR2_X1 i_4_0_222 (.A1(n_4_0_37), .A2(n_4_0_25), .ZN(\partial_reg[5] [24]));
   NOR2_X1 i_4_0_223 (.A1(n_4_0_37), .A2(n_4_0_26), .ZN(\partial_reg[5] [25]));
   NOR2_X1 i_4_0_224 (.A1(n_4_0_37), .A2(n_4_0_27), .ZN(\partial_reg[5] [26]));
   NOR2_X1 i_4_0_225 (.A1(n_4_0_37), .A2(n_4_0_28), .ZN(\partial_reg[5] [27]));
   NOR2_X1 i_4_0_226 (.A1(n_4_0_37), .A2(n_4_0_29), .ZN(\partial_reg[5] [28]));
   NOR2_X1 i_4_0_227 (.A1(n_4_0_37), .A2(n_4_0_30), .ZN(\partial_reg[5] [29]));
   NOR2_X1 i_4_0_228 (.A1(n_4_0_37), .A2(n_4_0_31), .ZN(\partial_reg[5] [30]));
   NOR2_X1 i_4_0_229 (.A1(n_4_0_37), .A2(n_4_0_32), .ZN(\partial_reg[5] [31]));
   INV_X1 i_4_0_230 (.A(op2[6]), .ZN(n_4_0_38));
   NOR2_X1 i_4_0_231 (.A1(n_4_0_38), .A2(n_4_0_1), .ZN(\partial_reg[6] [0]));
   NOR2_X1 i_4_0_232 (.A1(n_4_0_38), .A2(n_4_0_2), .ZN(\partial_reg[6] [1]));
   NOR2_X1 i_4_0_233 (.A1(n_4_0_38), .A2(n_4_0_3), .ZN(\partial_reg[6] [2]));
   NOR2_X1 i_4_0_234 (.A1(n_4_0_38), .A2(n_4_0_4), .ZN(\partial_reg[6] [3]));
   NOR2_X1 i_4_0_235 (.A1(n_4_0_38), .A2(n_4_0_5), .ZN(\partial_reg[6] [4]));
   NOR2_X1 i_4_0_236 (.A1(n_4_0_38), .A2(n_4_0_6), .ZN(\partial_reg[6] [5]));
   NOR2_X1 i_4_0_237 (.A1(n_4_0_38), .A2(n_4_0_7), .ZN(\partial_reg[6] [6]));
   NOR2_X1 i_4_0_238 (.A1(n_4_0_38), .A2(n_4_0_8), .ZN(\partial_reg[6] [7]));
   NOR2_X1 i_4_0_239 (.A1(n_4_0_38), .A2(n_4_0_9), .ZN(\partial_reg[6] [8]));
   NOR2_X1 i_4_0_240 (.A1(n_4_0_38), .A2(n_4_0_10), .ZN(\partial_reg[6] [9]));
   NOR2_X1 i_4_0_241 (.A1(n_4_0_38), .A2(n_4_0_11), .ZN(\partial_reg[6] [10]));
   NOR2_X1 i_4_0_242 (.A1(n_4_0_38), .A2(n_4_0_12), .ZN(\partial_reg[6] [11]));
   NOR2_X1 i_4_0_243 (.A1(n_4_0_38), .A2(n_4_0_13), .ZN(\partial_reg[6] [12]));
   NOR2_X1 i_4_0_244 (.A1(n_4_0_38), .A2(n_4_0_14), .ZN(\partial_reg[6] [13]));
   NOR2_X1 i_4_0_245 (.A1(n_4_0_38), .A2(n_4_0_15), .ZN(\partial_reg[6] [14]));
   NOR2_X1 i_4_0_246 (.A1(n_4_0_38), .A2(n_4_0_16), .ZN(\partial_reg[6] [15]));
   NOR2_X1 i_4_0_247 (.A1(n_4_0_38), .A2(n_4_0_17), .ZN(\partial_reg[6] [16]));
   NOR2_X1 i_4_0_248 (.A1(n_4_0_38), .A2(n_4_0_18), .ZN(\partial_reg[6] [17]));
   NOR2_X1 i_4_0_249 (.A1(n_4_0_38), .A2(n_4_0_19), .ZN(\partial_reg[6] [18]));
   NOR2_X1 i_4_0_250 (.A1(n_4_0_38), .A2(n_4_0_20), .ZN(\partial_reg[6] [19]));
   NOR2_X1 i_4_0_251 (.A1(n_4_0_38), .A2(n_4_0_21), .ZN(\partial_reg[6] [20]));
   NOR2_X1 i_4_0_252 (.A1(n_4_0_38), .A2(n_4_0_22), .ZN(\partial_reg[6] [21]));
   NOR2_X1 i_4_0_253 (.A1(n_4_0_38), .A2(n_4_0_23), .ZN(\partial_reg[6] [22]));
   NOR2_X1 i_4_0_254 (.A1(n_4_0_38), .A2(n_4_0_24), .ZN(\partial_reg[6] [23]));
   NOR2_X1 i_4_0_255 (.A1(n_4_0_38), .A2(n_4_0_25), .ZN(\partial_reg[6] [24]));
   NOR2_X1 i_4_0_256 (.A1(n_4_0_38), .A2(n_4_0_26), .ZN(\partial_reg[6] [25]));
   NOR2_X1 i_4_0_257 (.A1(n_4_0_38), .A2(n_4_0_27), .ZN(\partial_reg[6] [26]));
   NOR2_X1 i_4_0_258 (.A1(n_4_0_38), .A2(n_4_0_28), .ZN(\partial_reg[6] [27]));
   NOR2_X1 i_4_0_259 (.A1(n_4_0_38), .A2(n_4_0_29), .ZN(\partial_reg[6] [28]));
   NOR2_X1 i_4_0_260 (.A1(n_4_0_38), .A2(n_4_0_30), .ZN(\partial_reg[6] [29]));
   NOR2_X1 i_4_0_261 (.A1(n_4_0_38), .A2(n_4_0_31), .ZN(\partial_reg[6] [30]));
   NOR2_X1 i_4_0_262 (.A1(n_4_0_38), .A2(n_4_0_32), .ZN(\partial_reg[6] [31]));
   INV_X1 i_4_0_263 (.A(op2[7]), .ZN(n_4_0_39));
   NOR2_X1 i_4_0_264 (.A1(n_4_0_39), .A2(n_4_0_1), .ZN(\partial_reg[7] [0]));
   NOR2_X1 i_4_0_265 (.A1(n_4_0_39), .A2(n_4_0_2), .ZN(\partial_reg[7] [1]));
   NOR2_X1 i_4_0_266 (.A1(n_4_0_39), .A2(n_4_0_3), .ZN(\partial_reg[7] [2]));
   NOR2_X1 i_4_0_267 (.A1(n_4_0_39), .A2(n_4_0_4), .ZN(\partial_reg[7] [3]));
   NOR2_X1 i_4_0_268 (.A1(n_4_0_39), .A2(n_4_0_5), .ZN(\partial_reg[7] [4]));
   NOR2_X1 i_4_0_269 (.A1(n_4_0_39), .A2(n_4_0_6), .ZN(\partial_reg[7] [5]));
   NOR2_X1 i_4_0_270 (.A1(n_4_0_39), .A2(n_4_0_7), .ZN(\partial_reg[7] [6]));
   NOR2_X1 i_4_0_271 (.A1(n_4_0_39), .A2(n_4_0_8), .ZN(\partial_reg[7] [7]));
   NOR2_X1 i_4_0_272 (.A1(n_4_0_39), .A2(n_4_0_9), .ZN(\partial_reg[7] [8]));
   NOR2_X1 i_4_0_273 (.A1(n_4_0_39), .A2(n_4_0_10), .ZN(\partial_reg[7] [9]));
   NOR2_X1 i_4_0_274 (.A1(n_4_0_39), .A2(n_4_0_11), .ZN(\partial_reg[7] [10]));
   NOR2_X1 i_4_0_275 (.A1(n_4_0_39), .A2(n_4_0_12), .ZN(\partial_reg[7] [11]));
   NOR2_X1 i_4_0_276 (.A1(n_4_0_39), .A2(n_4_0_13), .ZN(\partial_reg[7] [12]));
   NOR2_X1 i_4_0_277 (.A1(n_4_0_39), .A2(n_4_0_14), .ZN(\partial_reg[7] [13]));
   NOR2_X1 i_4_0_278 (.A1(n_4_0_39), .A2(n_4_0_15), .ZN(\partial_reg[7] [14]));
   NOR2_X1 i_4_0_279 (.A1(n_4_0_39), .A2(n_4_0_16), .ZN(\partial_reg[7] [15]));
   NOR2_X1 i_4_0_280 (.A1(n_4_0_39), .A2(n_4_0_17), .ZN(\partial_reg[7] [16]));
   NOR2_X1 i_4_0_281 (.A1(n_4_0_39), .A2(n_4_0_18), .ZN(\partial_reg[7] [17]));
   NOR2_X1 i_4_0_282 (.A1(n_4_0_39), .A2(n_4_0_19), .ZN(\partial_reg[7] [18]));
   NOR2_X1 i_4_0_283 (.A1(n_4_0_39), .A2(n_4_0_20), .ZN(\partial_reg[7] [19]));
   NOR2_X1 i_4_0_284 (.A1(n_4_0_39), .A2(n_4_0_21), .ZN(\partial_reg[7] [20]));
   NOR2_X1 i_4_0_285 (.A1(n_4_0_39), .A2(n_4_0_22), .ZN(\partial_reg[7] [21]));
   NOR2_X1 i_4_0_286 (.A1(n_4_0_39), .A2(n_4_0_23), .ZN(\partial_reg[7] [22]));
   NOR2_X1 i_4_0_287 (.A1(n_4_0_39), .A2(n_4_0_24), .ZN(\partial_reg[7] [23]));
   NOR2_X1 i_4_0_288 (.A1(n_4_0_39), .A2(n_4_0_25), .ZN(\partial_reg[7] [24]));
   NOR2_X1 i_4_0_289 (.A1(n_4_0_39), .A2(n_4_0_26), .ZN(\partial_reg[7] [25]));
   NOR2_X1 i_4_0_290 (.A1(n_4_0_39), .A2(n_4_0_27), .ZN(\partial_reg[7] [26]));
   NOR2_X1 i_4_0_291 (.A1(n_4_0_39), .A2(n_4_0_28), .ZN(\partial_reg[7] [27]));
   NOR2_X1 i_4_0_292 (.A1(n_4_0_39), .A2(n_4_0_29), .ZN(\partial_reg[7] [28]));
   NOR2_X1 i_4_0_293 (.A1(n_4_0_39), .A2(n_4_0_30), .ZN(\partial_reg[7] [29]));
   NOR2_X1 i_4_0_294 (.A1(n_4_0_39), .A2(n_4_0_31), .ZN(\partial_reg[7] [30]));
   NOR2_X1 i_4_0_295 (.A1(n_4_0_39), .A2(n_4_0_32), .ZN(\partial_reg[7] [31]));
   INV_X1 i_4_0_296 (.A(op2[8]), .ZN(n_4_0_40));
   NOR2_X1 i_4_0_297 (.A1(n_4_0_40), .A2(n_4_0_1), .ZN(\partial_reg[8] [0]));
   NOR2_X1 i_4_0_298 (.A1(n_4_0_40), .A2(n_4_0_2), .ZN(\partial_reg[8] [1]));
   NOR2_X1 i_4_0_299 (.A1(n_4_0_40), .A2(n_4_0_3), .ZN(\partial_reg[8] [2]));
   NOR2_X1 i_4_0_300 (.A1(n_4_0_40), .A2(n_4_0_4), .ZN(\partial_reg[8] [3]));
   NOR2_X1 i_4_0_301 (.A1(n_4_0_40), .A2(n_4_0_5), .ZN(\partial_reg[8] [4]));
   NOR2_X1 i_4_0_302 (.A1(n_4_0_40), .A2(n_4_0_6), .ZN(\partial_reg[8] [5]));
   NOR2_X1 i_4_0_303 (.A1(n_4_0_40), .A2(n_4_0_7), .ZN(\partial_reg[8] [6]));
   NOR2_X1 i_4_0_304 (.A1(n_4_0_40), .A2(n_4_0_8), .ZN(\partial_reg[8] [7]));
   NOR2_X1 i_4_0_305 (.A1(n_4_0_40), .A2(n_4_0_9), .ZN(\partial_reg[8] [8]));
   NOR2_X1 i_4_0_306 (.A1(n_4_0_40), .A2(n_4_0_10), .ZN(\partial_reg[8] [9]));
   NOR2_X1 i_4_0_307 (.A1(n_4_0_40), .A2(n_4_0_11), .ZN(\partial_reg[8] [10]));
   NOR2_X1 i_4_0_308 (.A1(n_4_0_40), .A2(n_4_0_12), .ZN(\partial_reg[8] [11]));
   NOR2_X1 i_4_0_309 (.A1(n_4_0_40), .A2(n_4_0_13), .ZN(\partial_reg[8] [12]));
   NOR2_X1 i_4_0_310 (.A1(n_4_0_40), .A2(n_4_0_14), .ZN(\partial_reg[8] [13]));
   NOR2_X1 i_4_0_311 (.A1(n_4_0_40), .A2(n_4_0_15), .ZN(\partial_reg[8] [14]));
   NOR2_X1 i_4_0_312 (.A1(n_4_0_40), .A2(n_4_0_16), .ZN(\partial_reg[8] [15]));
   NOR2_X1 i_4_0_313 (.A1(n_4_0_40), .A2(n_4_0_17), .ZN(\partial_reg[8] [16]));
   NOR2_X1 i_4_0_314 (.A1(n_4_0_40), .A2(n_4_0_18), .ZN(\partial_reg[8] [17]));
   NOR2_X1 i_4_0_315 (.A1(n_4_0_40), .A2(n_4_0_19), .ZN(\partial_reg[8] [18]));
   NOR2_X1 i_4_0_316 (.A1(n_4_0_40), .A2(n_4_0_20), .ZN(\partial_reg[8] [19]));
   NOR2_X1 i_4_0_317 (.A1(n_4_0_40), .A2(n_4_0_21), .ZN(\partial_reg[8] [20]));
   NOR2_X1 i_4_0_318 (.A1(n_4_0_40), .A2(n_4_0_22), .ZN(\partial_reg[8] [21]));
   NOR2_X1 i_4_0_319 (.A1(n_4_0_40), .A2(n_4_0_23), .ZN(\partial_reg[8] [22]));
   NOR2_X1 i_4_0_320 (.A1(n_4_0_40), .A2(n_4_0_24), .ZN(\partial_reg[8] [23]));
   NOR2_X1 i_4_0_321 (.A1(n_4_0_40), .A2(n_4_0_25), .ZN(\partial_reg[8] [24]));
   NOR2_X1 i_4_0_322 (.A1(n_4_0_40), .A2(n_4_0_26), .ZN(\partial_reg[8] [25]));
   NOR2_X1 i_4_0_323 (.A1(n_4_0_40), .A2(n_4_0_27), .ZN(\partial_reg[8] [26]));
   NOR2_X1 i_4_0_324 (.A1(n_4_0_40), .A2(n_4_0_28), .ZN(\partial_reg[8] [27]));
   NOR2_X1 i_4_0_325 (.A1(n_4_0_40), .A2(n_4_0_29), .ZN(\partial_reg[8] [28]));
   NOR2_X1 i_4_0_326 (.A1(n_4_0_40), .A2(n_4_0_30), .ZN(\partial_reg[8] [29]));
   NOR2_X1 i_4_0_327 (.A1(n_4_0_40), .A2(n_4_0_31), .ZN(\partial_reg[8] [30]));
   NOR2_X1 i_4_0_328 (.A1(n_4_0_40), .A2(n_4_0_32), .ZN(\partial_reg[8] [31]));
   INV_X1 i_4_0_329 (.A(op2[9]), .ZN(n_4_0_41));
   NOR2_X1 i_4_0_330 (.A1(n_4_0_41), .A2(n_4_0_1), .ZN(\partial_reg[9] [0]));
   NOR2_X1 i_4_0_331 (.A1(n_4_0_41), .A2(n_4_0_2), .ZN(\partial_reg[9] [1]));
   NOR2_X1 i_4_0_332 (.A1(n_4_0_41), .A2(n_4_0_3), .ZN(\partial_reg[9] [2]));
   NOR2_X1 i_4_0_333 (.A1(n_4_0_41), .A2(n_4_0_4), .ZN(\partial_reg[9] [3]));
   NOR2_X1 i_4_0_334 (.A1(n_4_0_41), .A2(n_4_0_5), .ZN(\partial_reg[9] [4]));
   NOR2_X1 i_4_0_335 (.A1(n_4_0_41), .A2(n_4_0_6), .ZN(\partial_reg[9] [5]));
   NOR2_X1 i_4_0_336 (.A1(n_4_0_41), .A2(n_4_0_7), .ZN(\partial_reg[9] [6]));
   NOR2_X1 i_4_0_337 (.A1(n_4_0_41), .A2(n_4_0_8), .ZN(\partial_reg[9] [7]));
   NOR2_X1 i_4_0_338 (.A1(n_4_0_41), .A2(n_4_0_9), .ZN(\partial_reg[9] [8]));
   NOR2_X1 i_4_0_339 (.A1(n_4_0_41), .A2(n_4_0_10), .ZN(\partial_reg[9] [9]));
   NOR2_X1 i_4_0_340 (.A1(n_4_0_41), .A2(n_4_0_11), .ZN(\partial_reg[9] [10]));
   NOR2_X1 i_4_0_341 (.A1(n_4_0_41), .A2(n_4_0_12), .ZN(\partial_reg[9] [11]));
   NOR2_X1 i_4_0_342 (.A1(n_4_0_41), .A2(n_4_0_13), .ZN(\partial_reg[9] [12]));
   NOR2_X1 i_4_0_343 (.A1(n_4_0_41), .A2(n_4_0_14), .ZN(\partial_reg[9] [13]));
   NOR2_X1 i_4_0_344 (.A1(n_4_0_41), .A2(n_4_0_15), .ZN(\partial_reg[9] [14]));
   NOR2_X1 i_4_0_345 (.A1(n_4_0_41), .A2(n_4_0_16), .ZN(\partial_reg[9] [15]));
   NOR2_X1 i_4_0_346 (.A1(n_4_0_41), .A2(n_4_0_17), .ZN(\partial_reg[9] [16]));
   NOR2_X1 i_4_0_347 (.A1(n_4_0_41), .A2(n_4_0_18), .ZN(\partial_reg[9] [17]));
   NOR2_X1 i_4_0_348 (.A1(n_4_0_41), .A2(n_4_0_19), .ZN(\partial_reg[9] [18]));
   NOR2_X1 i_4_0_349 (.A1(n_4_0_41), .A2(n_4_0_20), .ZN(\partial_reg[9] [19]));
   NOR2_X1 i_4_0_350 (.A1(n_4_0_41), .A2(n_4_0_21), .ZN(\partial_reg[9] [20]));
   NOR2_X1 i_4_0_351 (.A1(n_4_0_41), .A2(n_4_0_22), .ZN(\partial_reg[9] [21]));
   NOR2_X1 i_4_0_352 (.A1(n_4_0_41), .A2(n_4_0_23), .ZN(\partial_reg[9] [22]));
   NOR2_X1 i_4_0_353 (.A1(n_4_0_41), .A2(n_4_0_24), .ZN(\partial_reg[9] [23]));
   NOR2_X1 i_4_0_354 (.A1(n_4_0_41), .A2(n_4_0_25), .ZN(\partial_reg[9] [24]));
   NOR2_X1 i_4_0_355 (.A1(n_4_0_41), .A2(n_4_0_26), .ZN(\partial_reg[9] [25]));
   NOR2_X1 i_4_0_356 (.A1(n_4_0_41), .A2(n_4_0_27), .ZN(\partial_reg[9] [26]));
   NOR2_X1 i_4_0_357 (.A1(n_4_0_41), .A2(n_4_0_28), .ZN(\partial_reg[9] [27]));
   NOR2_X1 i_4_0_358 (.A1(n_4_0_41), .A2(n_4_0_29), .ZN(\partial_reg[9] [28]));
   NOR2_X1 i_4_0_359 (.A1(n_4_0_41), .A2(n_4_0_30), .ZN(\partial_reg[9] [29]));
   NOR2_X1 i_4_0_360 (.A1(n_4_0_41), .A2(n_4_0_31), .ZN(\partial_reg[9] [30]));
   NOR2_X1 i_4_0_361 (.A1(n_4_0_41), .A2(n_4_0_32), .ZN(\partial_reg[9] [31]));
   INV_X1 i_4_0_362 (.A(op2[10]), .ZN(n_4_0_42));
   NOR2_X1 i_4_0_363 (.A1(n_4_0_42), .A2(n_4_0_1), .ZN(\partial_reg[10] [0]));
   NOR2_X1 i_4_0_364 (.A1(n_4_0_42), .A2(n_4_0_2), .ZN(\partial_reg[10] [1]));
   NOR2_X1 i_4_0_365 (.A1(n_4_0_42), .A2(n_4_0_3), .ZN(\partial_reg[10] [2]));
   NOR2_X1 i_4_0_366 (.A1(n_4_0_42), .A2(n_4_0_4), .ZN(\partial_reg[10] [3]));
   NOR2_X1 i_4_0_367 (.A1(n_4_0_42), .A2(n_4_0_5), .ZN(\partial_reg[10] [4]));
   NOR2_X1 i_4_0_368 (.A1(n_4_0_42), .A2(n_4_0_6), .ZN(\partial_reg[10] [5]));
   NOR2_X1 i_4_0_369 (.A1(n_4_0_42), .A2(n_4_0_7), .ZN(\partial_reg[10] [6]));
   NOR2_X1 i_4_0_370 (.A1(n_4_0_42), .A2(n_4_0_8), .ZN(\partial_reg[10] [7]));
   NOR2_X1 i_4_0_371 (.A1(n_4_0_42), .A2(n_4_0_9), .ZN(\partial_reg[10] [8]));
   NOR2_X1 i_4_0_372 (.A1(n_4_0_42), .A2(n_4_0_10), .ZN(\partial_reg[10] [9]));
   NOR2_X1 i_4_0_373 (.A1(n_4_0_42), .A2(n_4_0_11), .ZN(\partial_reg[10] [10]));
   NOR2_X1 i_4_0_374 (.A1(n_4_0_42), .A2(n_4_0_12), .ZN(\partial_reg[10] [11]));
   NOR2_X1 i_4_0_375 (.A1(n_4_0_42), .A2(n_4_0_13), .ZN(\partial_reg[10] [12]));
   NOR2_X1 i_4_0_376 (.A1(n_4_0_42), .A2(n_4_0_14), .ZN(\partial_reg[10] [13]));
   NOR2_X1 i_4_0_377 (.A1(n_4_0_42), .A2(n_4_0_15), .ZN(\partial_reg[10] [14]));
   NOR2_X1 i_4_0_378 (.A1(n_4_0_42), .A2(n_4_0_16), .ZN(\partial_reg[10] [15]));
   NOR2_X1 i_4_0_379 (.A1(n_4_0_42), .A2(n_4_0_17), .ZN(\partial_reg[10] [16]));
   NOR2_X1 i_4_0_380 (.A1(n_4_0_42), .A2(n_4_0_18), .ZN(\partial_reg[10] [17]));
   NOR2_X1 i_4_0_381 (.A1(n_4_0_42), .A2(n_4_0_19), .ZN(\partial_reg[10] [18]));
   NOR2_X1 i_4_0_382 (.A1(n_4_0_42), .A2(n_4_0_20), .ZN(\partial_reg[10] [19]));
   NOR2_X1 i_4_0_383 (.A1(n_4_0_42), .A2(n_4_0_21), .ZN(\partial_reg[10] [20]));
   NOR2_X1 i_4_0_384 (.A1(n_4_0_42), .A2(n_4_0_22), .ZN(\partial_reg[10] [21]));
   NOR2_X1 i_4_0_385 (.A1(n_4_0_42), .A2(n_4_0_23), .ZN(\partial_reg[10] [22]));
   NOR2_X1 i_4_0_386 (.A1(n_4_0_42), .A2(n_4_0_24), .ZN(\partial_reg[10] [23]));
   NOR2_X1 i_4_0_387 (.A1(n_4_0_42), .A2(n_4_0_25), .ZN(\partial_reg[10] [24]));
   NOR2_X1 i_4_0_388 (.A1(n_4_0_42), .A2(n_4_0_26), .ZN(\partial_reg[10] [25]));
   NOR2_X1 i_4_0_389 (.A1(n_4_0_42), .A2(n_4_0_27), .ZN(\partial_reg[10] [26]));
   NOR2_X1 i_4_0_390 (.A1(n_4_0_42), .A2(n_4_0_28), .ZN(\partial_reg[10] [27]));
   NOR2_X1 i_4_0_391 (.A1(n_4_0_42), .A2(n_4_0_29), .ZN(\partial_reg[10] [28]));
   NOR2_X1 i_4_0_392 (.A1(n_4_0_42), .A2(n_4_0_30), .ZN(\partial_reg[10] [29]));
   NOR2_X1 i_4_0_393 (.A1(n_4_0_42), .A2(n_4_0_31), .ZN(\partial_reg[10] [30]));
   NOR2_X1 i_4_0_394 (.A1(n_4_0_42), .A2(n_4_0_32), .ZN(\partial_reg[10] [31]));
   INV_X1 i_4_0_395 (.A(op2[11]), .ZN(n_4_0_43));
   NOR2_X1 i_4_0_396 (.A1(n_4_0_43), .A2(n_4_0_1), .ZN(\partial_reg[11] [0]));
   NOR2_X1 i_4_0_397 (.A1(n_4_0_43), .A2(n_4_0_2), .ZN(\partial_reg[11] [1]));
   NOR2_X1 i_4_0_398 (.A1(n_4_0_43), .A2(n_4_0_3), .ZN(\partial_reg[11] [2]));
   NOR2_X1 i_4_0_399 (.A1(n_4_0_43), .A2(n_4_0_4), .ZN(\partial_reg[11] [3]));
   NOR2_X1 i_4_0_400 (.A1(n_4_0_43), .A2(n_4_0_5), .ZN(\partial_reg[11] [4]));
   NOR2_X1 i_4_0_401 (.A1(n_4_0_43), .A2(n_4_0_6), .ZN(\partial_reg[11] [5]));
   NOR2_X1 i_4_0_402 (.A1(n_4_0_43), .A2(n_4_0_7), .ZN(\partial_reg[11] [6]));
   NOR2_X1 i_4_0_403 (.A1(n_4_0_43), .A2(n_4_0_8), .ZN(\partial_reg[11] [7]));
   NOR2_X1 i_4_0_404 (.A1(n_4_0_43), .A2(n_4_0_9), .ZN(\partial_reg[11] [8]));
   NOR2_X1 i_4_0_405 (.A1(n_4_0_43), .A2(n_4_0_10), .ZN(\partial_reg[11] [9]));
   NOR2_X1 i_4_0_406 (.A1(n_4_0_43), .A2(n_4_0_11), .ZN(\partial_reg[11] [10]));
   NOR2_X1 i_4_0_407 (.A1(n_4_0_43), .A2(n_4_0_12), .ZN(\partial_reg[11] [11]));
   NOR2_X1 i_4_0_408 (.A1(n_4_0_43), .A2(n_4_0_13), .ZN(\partial_reg[11] [12]));
   NOR2_X1 i_4_0_409 (.A1(n_4_0_43), .A2(n_4_0_14), .ZN(\partial_reg[11] [13]));
   NOR2_X1 i_4_0_410 (.A1(n_4_0_43), .A2(n_4_0_15), .ZN(\partial_reg[11] [14]));
   NOR2_X1 i_4_0_411 (.A1(n_4_0_43), .A2(n_4_0_16), .ZN(\partial_reg[11] [15]));
   NOR2_X1 i_4_0_412 (.A1(n_4_0_43), .A2(n_4_0_17), .ZN(\partial_reg[11] [16]));
   NOR2_X1 i_4_0_413 (.A1(n_4_0_43), .A2(n_4_0_18), .ZN(\partial_reg[11] [17]));
   NOR2_X1 i_4_0_414 (.A1(n_4_0_43), .A2(n_4_0_19), .ZN(\partial_reg[11] [18]));
   NOR2_X1 i_4_0_415 (.A1(n_4_0_43), .A2(n_4_0_20), .ZN(\partial_reg[11] [19]));
   NOR2_X1 i_4_0_416 (.A1(n_4_0_43), .A2(n_4_0_21), .ZN(\partial_reg[11] [20]));
   NOR2_X1 i_4_0_417 (.A1(n_4_0_43), .A2(n_4_0_22), .ZN(\partial_reg[11] [21]));
   NOR2_X1 i_4_0_418 (.A1(n_4_0_43), .A2(n_4_0_23), .ZN(\partial_reg[11] [22]));
   NOR2_X1 i_4_0_419 (.A1(n_4_0_43), .A2(n_4_0_24), .ZN(\partial_reg[11] [23]));
   NOR2_X1 i_4_0_420 (.A1(n_4_0_43), .A2(n_4_0_25), .ZN(\partial_reg[11] [24]));
   NOR2_X1 i_4_0_421 (.A1(n_4_0_43), .A2(n_4_0_26), .ZN(\partial_reg[11] [25]));
   NOR2_X1 i_4_0_422 (.A1(n_4_0_43), .A2(n_4_0_27), .ZN(\partial_reg[11] [26]));
   NOR2_X1 i_4_0_423 (.A1(n_4_0_43), .A2(n_4_0_28), .ZN(\partial_reg[11] [27]));
   NOR2_X1 i_4_0_424 (.A1(n_4_0_43), .A2(n_4_0_29), .ZN(\partial_reg[11] [28]));
   NOR2_X1 i_4_0_425 (.A1(n_4_0_43), .A2(n_4_0_30), .ZN(\partial_reg[11] [29]));
   NOR2_X1 i_4_0_426 (.A1(n_4_0_43), .A2(n_4_0_31), .ZN(\partial_reg[11] [30]));
   NOR2_X1 i_4_0_427 (.A1(n_4_0_43), .A2(n_4_0_32), .ZN(\partial_reg[11] [31]));
   INV_X1 i_4_0_428 (.A(op2[12]), .ZN(n_4_0_44));
   NOR2_X1 i_4_0_429 (.A1(n_4_0_44), .A2(n_4_0_1), .ZN(\partial_reg[12] [0]));
   NOR2_X1 i_4_0_430 (.A1(n_4_0_44), .A2(n_4_0_2), .ZN(\partial_reg[12] [1]));
   NOR2_X1 i_4_0_431 (.A1(n_4_0_44), .A2(n_4_0_3), .ZN(\partial_reg[12] [2]));
   NOR2_X1 i_4_0_432 (.A1(n_4_0_44), .A2(n_4_0_4), .ZN(\partial_reg[12] [3]));
   NOR2_X1 i_4_0_433 (.A1(n_4_0_44), .A2(n_4_0_5), .ZN(\partial_reg[12] [4]));
   NOR2_X1 i_4_0_434 (.A1(n_4_0_44), .A2(n_4_0_6), .ZN(\partial_reg[12] [5]));
   NOR2_X1 i_4_0_435 (.A1(n_4_0_44), .A2(n_4_0_7), .ZN(\partial_reg[12] [6]));
   NOR2_X1 i_4_0_436 (.A1(n_4_0_44), .A2(n_4_0_8), .ZN(\partial_reg[12] [7]));
   NOR2_X1 i_4_0_437 (.A1(n_4_0_44), .A2(n_4_0_9), .ZN(\partial_reg[12] [8]));
   NOR2_X1 i_4_0_438 (.A1(n_4_0_44), .A2(n_4_0_10), .ZN(\partial_reg[12] [9]));
   NOR2_X1 i_4_0_439 (.A1(n_4_0_44), .A2(n_4_0_11), .ZN(\partial_reg[12] [10]));
   NOR2_X1 i_4_0_440 (.A1(n_4_0_44), .A2(n_4_0_12), .ZN(\partial_reg[12] [11]));
   NOR2_X1 i_4_0_441 (.A1(n_4_0_44), .A2(n_4_0_13), .ZN(\partial_reg[12] [12]));
   NOR2_X1 i_4_0_442 (.A1(n_4_0_44), .A2(n_4_0_14), .ZN(\partial_reg[12] [13]));
   NOR2_X1 i_4_0_443 (.A1(n_4_0_44), .A2(n_4_0_15), .ZN(\partial_reg[12] [14]));
   NOR2_X1 i_4_0_444 (.A1(n_4_0_44), .A2(n_4_0_16), .ZN(\partial_reg[12] [15]));
   NOR2_X1 i_4_0_445 (.A1(n_4_0_44), .A2(n_4_0_17), .ZN(\partial_reg[12] [16]));
   NOR2_X1 i_4_0_446 (.A1(n_4_0_44), .A2(n_4_0_18), .ZN(\partial_reg[12] [17]));
   NOR2_X1 i_4_0_447 (.A1(n_4_0_44), .A2(n_4_0_19), .ZN(\partial_reg[12] [18]));
   NOR2_X1 i_4_0_448 (.A1(n_4_0_44), .A2(n_4_0_20), .ZN(\partial_reg[12] [19]));
   NOR2_X1 i_4_0_449 (.A1(n_4_0_44), .A2(n_4_0_21), .ZN(\partial_reg[12] [20]));
   NOR2_X1 i_4_0_450 (.A1(n_4_0_44), .A2(n_4_0_22), .ZN(\partial_reg[12] [21]));
   NOR2_X1 i_4_0_451 (.A1(n_4_0_44), .A2(n_4_0_23), .ZN(\partial_reg[12] [22]));
   NOR2_X1 i_4_0_452 (.A1(n_4_0_44), .A2(n_4_0_24), .ZN(\partial_reg[12] [23]));
   NOR2_X1 i_4_0_453 (.A1(n_4_0_44), .A2(n_4_0_25), .ZN(\partial_reg[12] [24]));
   NOR2_X1 i_4_0_454 (.A1(n_4_0_44), .A2(n_4_0_26), .ZN(\partial_reg[12] [25]));
   NOR2_X1 i_4_0_455 (.A1(n_4_0_44), .A2(n_4_0_27), .ZN(\partial_reg[12] [26]));
   NOR2_X1 i_4_0_456 (.A1(n_4_0_44), .A2(n_4_0_28), .ZN(\partial_reg[12] [27]));
   NOR2_X1 i_4_0_457 (.A1(n_4_0_44), .A2(n_4_0_29), .ZN(\partial_reg[12] [28]));
   NOR2_X1 i_4_0_458 (.A1(n_4_0_44), .A2(n_4_0_30), .ZN(\partial_reg[12] [29]));
   NOR2_X1 i_4_0_459 (.A1(n_4_0_44), .A2(n_4_0_31), .ZN(\partial_reg[12] [30]));
   NOR2_X1 i_4_0_460 (.A1(n_4_0_44), .A2(n_4_0_32), .ZN(\partial_reg[12] [31]));
   INV_X1 i_4_0_461 (.A(op2[13]), .ZN(n_4_0_45));
   NOR2_X1 i_4_0_462 (.A1(n_4_0_45), .A2(n_4_0_1), .ZN(\partial_reg[13] [0]));
   NOR2_X1 i_4_0_463 (.A1(n_4_0_45), .A2(n_4_0_2), .ZN(\partial_reg[13] [1]));
   NOR2_X1 i_4_0_464 (.A1(n_4_0_45), .A2(n_4_0_3), .ZN(\partial_reg[13] [2]));
   NOR2_X1 i_4_0_465 (.A1(n_4_0_45), .A2(n_4_0_4), .ZN(\partial_reg[13] [3]));
   NOR2_X1 i_4_0_466 (.A1(n_4_0_45), .A2(n_4_0_5), .ZN(\partial_reg[13] [4]));
   NOR2_X1 i_4_0_467 (.A1(n_4_0_45), .A2(n_4_0_6), .ZN(\partial_reg[13] [5]));
   NOR2_X1 i_4_0_468 (.A1(n_4_0_45), .A2(n_4_0_7), .ZN(\partial_reg[13] [6]));
   NOR2_X1 i_4_0_469 (.A1(n_4_0_45), .A2(n_4_0_8), .ZN(\partial_reg[13] [7]));
   NOR2_X1 i_4_0_470 (.A1(n_4_0_45), .A2(n_4_0_9), .ZN(\partial_reg[13] [8]));
   NOR2_X1 i_4_0_471 (.A1(n_4_0_45), .A2(n_4_0_10), .ZN(\partial_reg[13] [9]));
   NOR2_X1 i_4_0_472 (.A1(n_4_0_45), .A2(n_4_0_11), .ZN(\partial_reg[13] [10]));
   NOR2_X1 i_4_0_473 (.A1(n_4_0_45), .A2(n_4_0_12), .ZN(\partial_reg[13] [11]));
   NOR2_X1 i_4_0_474 (.A1(n_4_0_45), .A2(n_4_0_13), .ZN(\partial_reg[13] [12]));
   NOR2_X1 i_4_0_475 (.A1(n_4_0_45), .A2(n_4_0_14), .ZN(\partial_reg[13] [13]));
   NOR2_X1 i_4_0_476 (.A1(n_4_0_45), .A2(n_4_0_15), .ZN(\partial_reg[13] [14]));
   NOR2_X1 i_4_0_477 (.A1(n_4_0_45), .A2(n_4_0_16), .ZN(\partial_reg[13] [15]));
   NOR2_X1 i_4_0_478 (.A1(n_4_0_45), .A2(n_4_0_17), .ZN(\partial_reg[13] [16]));
   NOR2_X1 i_4_0_479 (.A1(n_4_0_45), .A2(n_4_0_18), .ZN(\partial_reg[13] [17]));
   NOR2_X1 i_4_0_480 (.A1(n_4_0_45), .A2(n_4_0_19), .ZN(\partial_reg[13] [18]));
   NOR2_X1 i_4_0_481 (.A1(n_4_0_45), .A2(n_4_0_20), .ZN(\partial_reg[13] [19]));
   NOR2_X1 i_4_0_482 (.A1(n_4_0_45), .A2(n_4_0_21), .ZN(\partial_reg[13] [20]));
   NOR2_X1 i_4_0_483 (.A1(n_4_0_45), .A2(n_4_0_22), .ZN(\partial_reg[13] [21]));
   NOR2_X1 i_4_0_484 (.A1(n_4_0_45), .A2(n_4_0_23), .ZN(\partial_reg[13] [22]));
   NOR2_X1 i_4_0_485 (.A1(n_4_0_45), .A2(n_4_0_24), .ZN(\partial_reg[13] [23]));
   NOR2_X1 i_4_0_486 (.A1(n_4_0_45), .A2(n_4_0_25), .ZN(\partial_reg[13] [24]));
   NOR2_X1 i_4_0_487 (.A1(n_4_0_45), .A2(n_4_0_26), .ZN(\partial_reg[13] [25]));
   NOR2_X1 i_4_0_488 (.A1(n_4_0_45), .A2(n_4_0_27), .ZN(\partial_reg[13] [26]));
   NOR2_X1 i_4_0_489 (.A1(n_4_0_45), .A2(n_4_0_28), .ZN(\partial_reg[13] [27]));
   NOR2_X1 i_4_0_490 (.A1(n_4_0_45), .A2(n_4_0_29), .ZN(\partial_reg[13] [28]));
   NOR2_X1 i_4_0_491 (.A1(n_4_0_45), .A2(n_4_0_30), .ZN(\partial_reg[13] [29]));
   NOR2_X1 i_4_0_492 (.A1(n_4_0_45), .A2(n_4_0_31), .ZN(\partial_reg[13] [30]));
   NOR2_X1 i_4_0_493 (.A1(n_4_0_45), .A2(n_4_0_32), .ZN(\partial_reg[13] [31]));
   INV_X1 i_4_0_494 (.A(op2[14]), .ZN(n_4_0_46));
   NOR2_X1 i_4_0_495 (.A1(n_4_0_46), .A2(n_4_0_1), .ZN(\partial_reg[14] [0]));
   NOR2_X1 i_4_0_496 (.A1(n_4_0_46), .A2(n_4_0_2), .ZN(\partial_reg[14] [1]));
   NOR2_X1 i_4_0_497 (.A1(n_4_0_46), .A2(n_4_0_3), .ZN(\partial_reg[14] [2]));
   NOR2_X1 i_4_0_498 (.A1(n_4_0_46), .A2(n_4_0_4), .ZN(\partial_reg[14] [3]));
   NOR2_X1 i_4_0_499 (.A1(n_4_0_46), .A2(n_4_0_5), .ZN(\partial_reg[14] [4]));
   NOR2_X1 i_4_0_500 (.A1(n_4_0_46), .A2(n_4_0_6), .ZN(\partial_reg[14] [5]));
   NOR2_X1 i_4_0_501 (.A1(n_4_0_46), .A2(n_4_0_7), .ZN(\partial_reg[14] [6]));
   NOR2_X1 i_4_0_502 (.A1(n_4_0_46), .A2(n_4_0_8), .ZN(\partial_reg[14] [7]));
   NOR2_X1 i_4_0_503 (.A1(n_4_0_46), .A2(n_4_0_9), .ZN(\partial_reg[14] [8]));
   NOR2_X1 i_4_0_504 (.A1(n_4_0_46), .A2(n_4_0_10), .ZN(\partial_reg[14] [9]));
   NOR2_X1 i_4_0_505 (.A1(n_4_0_46), .A2(n_4_0_11), .ZN(\partial_reg[14] [10]));
   NOR2_X1 i_4_0_506 (.A1(n_4_0_46), .A2(n_4_0_12), .ZN(\partial_reg[14] [11]));
   NOR2_X1 i_4_0_507 (.A1(n_4_0_46), .A2(n_4_0_13), .ZN(\partial_reg[14] [12]));
   NOR2_X1 i_4_0_508 (.A1(n_4_0_46), .A2(n_4_0_14), .ZN(\partial_reg[14] [13]));
   NOR2_X1 i_4_0_509 (.A1(n_4_0_46), .A2(n_4_0_15), .ZN(\partial_reg[14] [14]));
   NOR2_X1 i_4_0_510 (.A1(n_4_0_46), .A2(n_4_0_16), .ZN(\partial_reg[14] [15]));
   NOR2_X1 i_4_0_511 (.A1(n_4_0_46), .A2(n_4_0_17), .ZN(\partial_reg[14] [16]));
   NOR2_X1 i_4_0_512 (.A1(n_4_0_46), .A2(n_4_0_18), .ZN(\partial_reg[14] [17]));
   NOR2_X1 i_4_0_513 (.A1(n_4_0_46), .A2(n_4_0_19), .ZN(\partial_reg[14] [18]));
   NOR2_X1 i_4_0_514 (.A1(n_4_0_46), .A2(n_4_0_20), .ZN(\partial_reg[14] [19]));
   NOR2_X1 i_4_0_515 (.A1(n_4_0_46), .A2(n_4_0_21), .ZN(\partial_reg[14] [20]));
   NOR2_X1 i_4_0_516 (.A1(n_4_0_46), .A2(n_4_0_22), .ZN(\partial_reg[14] [21]));
   NOR2_X1 i_4_0_517 (.A1(n_4_0_46), .A2(n_4_0_23), .ZN(\partial_reg[14] [22]));
   NOR2_X1 i_4_0_518 (.A1(n_4_0_46), .A2(n_4_0_24), .ZN(\partial_reg[14] [23]));
   NOR2_X1 i_4_0_519 (.A1(n_4_0_46), .A2(n_4_0_25), .ZN(\partial_reg[14] [24]));
   NOR2_X1 i_4_0_520 (.A1(n_4_0_46), .A2(n_4_0_26), .ZN(\partial_reg[14] [25]));
   NOR2_X1 i_4_0_521 (.A1(n_4_0_46), .A2(n_4_0_27), .ZN(\partial_reg[14] [26]));
   NOR2_X1 i_4_0_522 (.A1(n_4_0_46), .A2(n_4_0_28), .ZN(\partial_reg[14] [27]));
   NOR2_X1 i_4_0_523 (.A1(n_4_0_46), .A2(n_4_0_29), .ZN(\partial_reg[14] [28]));
   NOR2_X1 i_4_0_524 (.A1(n_4_0_46), .A2(n_4_0_30), .ZN(\partial_reg[14] [29]));
   NOR2_X1 i_4_0_525 (.A1(n_4_0_46), .A2(n_4_0_31), .ZN(\partial_reg[14] [30]));
   NOR2_X1 i_4_0_526 (.A1(n_4_0_46), .A2(n_4_0_32), .ZN(\partial_reg[14] [31]));
   INV_X1 i_4_0_527 (.A(op2[15]), .ZN(n_4_0_47));
   NOR2_X1 i_4_0_528 (.A1(n_4_0_47), .A2(n_4_0_1), .ZN(\partial_reg[15] [0]));
   NOR2_X1 i_4_0_529 (.A1(n_4_0_47), .A2(n_4_0_2), .ZN(\partial_reg[15] [1]));
   NOR2_X1 i_4_0_530 (.A1(n_4_0_47), .A2(n_4_0_3), .ZN(\partial_reg[15] [2]));
   NOR2_X1 i_4_0_531 (.A1(n_4_0_47), .A2(n_4_0_4), .ZN(\partial_reg[15] [3]));
   NOR2_X1 i_4_0_532 (.A1(n_4_0_47), .A2(n_4_0_5), .ZN(\partial_reg[15] [4]));
   NOR2_X1 i_4_0_533 (.A1(n_4_0_47), .A2(n_4_0_6), .ZN(\partial_reg[15] [5]));
   NOR2_X1 i_4_0_534 (.A1(n_4_0_47), .A2(n_4_0_7), .ZN(\partial_reg[15] [6]));
   NOR2_X1 i_4_0_535 (.A1(n_4_0_47), .A2(n_4_0_8), .ZN(\partial_reg[15] [7]));
   NOR2_X1 i_4_0_536 (.A1(n_4_0_47), .A2(n_4_0_9), .ZN(\partial_reg[15] [8]));
   NOR2_X1 i_4_0_537 (.A1(n_4_0_47), .A2(n_4_0_10), .ZN(\partial_reg[15] [9]));
   NOR2_X1 i_4_0_538 (.A1(n_4_0_47), .A2(n_4_0_11), .ZN(\partial_reg[15] [10]));
   NOR2_X1 i_4_0_539 (.A1(n_4_0_47), .A2(n_4_0_12), .ZN(\partial_reg[15] [11]));
   NOR2_X1 i_4_0_540 (.A1(n_4_0_47), .A2(n_4_0_13), .ZN(\partial_reg[15] [12]));
   NOR2_X1 i_4_0_541 (.A1(n_4_0_47), .A2(n_4_0_14), .ZN(\partial_reg[15] [13]));
   NOR2_X1 i_4_0_542 (.A1(n_4_0_47), .A2(n_4_0_15), .ZN(\partial_reg[15] [14]));
   NOR2_X1 i_4_0_543 (.A1(n_4_0_47), .A2(n_4_0_16), .ZN(\partial_reg[15] [15]));
   NOR2_X1 i_4_0_544 (.A1(n_4_0_47), .A2(n_4_0_17), .ZN(\partial_reg[15] [16]));
   NOR2_X1 i_4_0_545 (.A1(n_4_0_47), .A2(n_4_0_18), .ZN(\partial_reg[15] [17]));
   NOR2_X1 i_4_0_546 (.A1(n_4_0_47), .A2(n_4_0_19), .ZN(\partial_reg[15] [18]));
   NOR2_X1 i_4_0_547 (.A1(n_4_0_47), .A2(n_4_0_20), .ZN(\partial_reg[15] [19]));
   NOR2_X1 i_4_0_548 (.A1(n_4_0_47), .A2(n_4_0_21), .ZN(\partial_reg[15] [20]));
   NOR2_X1 i_4_0_549 (.A1(n_4_0_47), .A2(n_4_0_22), .ZN(\partial_reg[15] [21]));
   NOR2_X1 i_4_0_550 (.A1(n_4_0_47), .A2(n_4_0_23), .ZN(\partial_reg[15] [22]));
   NOR2_X1 i_4_0_551 (.A1(n_4_0_47), .A2(n_4_0_24), .ZN(\partial_reg[15] [23]));
   NOR2_X1 i_4_0_552 (.A1(n_4_0_47), .A2(n_4_0_25), .ZN(\partial_reg[15] [24]));
   NOR2_X1 i_4_0_553 (.A1(n_4_0_47), .A2(n_4_0_26), .ZN(\partial_reg[15] [25]));
   NOR2_X1 i_4_0_554 (.A1(n_4_0_47), .A2(n_4_0_27), .ZN(\partial_reg[15] [26]));
   NOR2_X1 i_4_0_555 (.A1(n_4_0_47), .A2(n_4_0_28), .ZN(\partial_reg[15] [27]));
   NOR2_X1 i_4_0_556 (.A1(n_4_0_47), .A2(n_4_0_29), .ZN(\partial_reg[15] [28]));
   NOR2_X1 i_4_0_557 (.A1(n_4_0_47), .A2(n_4_0_30), .ZN(\partial_reg[15] [29]));
   NOR2_X1 i_4_0_558 (.A1(n_4_0_47), .A2(n_4_0_31), .ZN(\partial_reg[15] [30]));
   NOR2_X1 i_4_0_559 (.A1(n_4_0_47), .A2(n_4_0_32), .ZN(\partial_reg[15] [31]));
   INV_X1 i_4_0_560 (.A(op2[16]), .ZN(n_4_0_48));
   NOR2_X1 i_4_0_561 (.A1(n_4_0_48), .A2(n_4_0_1), .ZN(\partial_reg[16] [0]));
   NOR2_X1 i_4_0_562 (.A1(n_4_0_48), .A2(n_4_0_2), .ZN(\partial_reg[16] [1]));
   NOR2_X1 i_4_0_563 (.A1(n_4_0_48), .A2(n_4_0_3), .ZN(\partial_reg[16] [2]));
   NOR2_X1 i_4_0_564 (.A1(n_4_0_48), .A2(n_4_0_4), .ZN(\partial_reg[16] [3]));
   NOR2_X1 i_4_0_565 (.A1(n_4_0_48), .A2(n_4_0_5), .ZN(\partial_reg[16] [4]));
   NOR2_X1 i_4_0_566 (.A1(n_4_0_48), .A2(n_4_0_6), .ZN(\partial_reg[16] [5]));
   NOR2_X1 i_4_0_567 (.A1(n_4_0_48), .A2(n_4_0_7), .ZN(\partial_reg[16] [6]));
   NOR2_X1 i_4_0_568 (.A1(n_4_0_48), .A2(n_4_0_8), .ZN(\partial_reg[16] [7]));
   NOR2_X1 i_4_0_569 (.A1(n_4_0_48), .A2(n_4_0_9), .ZN(\partial_reg[16] [8]));
   NOR2_X1 i_4_0_570 (.A1(n_4_0_48), .A2(n_4_0_10), .ZN(\partial_reg[16] [9]));
   NOR2_X1 i_4_0_571 (.A1(n_4_0_48), .A2(n_4_0_11), .ZN(\partial_reg[16] [10]));
   NOR2_X1 i_4_0_572 (.A1(n_4_0_48), .A2(n_4_0_12), .ZN(\partial_reg[16] [11]));
   NOR2_X1 i_4_0_573 (.A1(n_4_0_48), .A2(n_4_0_13), .ZN(\partial_reg[16] [12]));
   NOR2_X1 i_4_0_574 (.A1(n_4_0_48), .A2(n_4_0_14), .ZN(\partial_reg[16] [13]));
   NOR2_X1 i_4_0_575 (.A1(n_4_0_48), .A2(n_4_0_15), .ZN(\partial_reg[16] [14]));
   NOR2_X1 i_4_0_576 (.A1(n_4_0_48), .A2(n_4_0_16), .ZN(\partial_reg[16] [15]));
   NOR2_X1 i_4_0_577 (.A1(n_4_0_48), .A2(n_4_0_17), .ZN(\partial_reg[16] [16]));
   NOR2_X1 i_4_0_578 (.A1(n_4_0_48), .A2(n_4_0_18), .ZN(\partial_reg[16] [17]));
   NOR2_X1 i_4_0_579 (.A1(n_4_0_48), .A2(n_4_0_19), .ZN(\partial_reg[16] [18]));
   NOR2_X1 i_4_0_580 (.A1(n_4_0_48), .A2(n_4_0_20), .ZN(\partial_reg[16] [19]));
   NOR2_X1 i_4_0_581 (.A1(n_4_0_48), .A2(n_4_0_21), .ZN(\partial_reg[16] [20]));
   NOR2_X1 i_4_0_582 (.A1(n_4_0_48), .A2(n_4_0_22), .ZN(\partial_reg[16] [21]));
   NOR2_X1 i_4_0_583 (.A1(n_4_0_48), .A2(n_4_0_23), .ZN(\partial_reg[16] [22]));
   NOR2_X1 i_4_0_584 (.A1(n_4_0_48), .A2(n_4_0_24), .ZN(\partial_reg[16] [23]));
   NOR2_X1 i_4_0_585 (.A1(n_4_0_48), .A2(n_4_0_25), .ZN(\partial_reg[16] [24]));
   NOR2_X1 i_4_0_586 (.A1(n_4_0_48), .A2(n_4_0_26), .ZN(\partial_reg[16] [25]));
   NOR2_X1 i_4_0_587 (.A1(n_4_0_48), .A2(n_4_0_27), .ZN(\partial_reg[16] [26]));
   NOR2_X1 i_4_0_588 (.A1(n_4_0_48), .A2(n_4_0_28), .ZN(\partial_reg[16] [27]));
   NOR2_X1 i_4_0_589 (.A1(n_4_0_48), .A2(n_4_0_29), .ZN(\partial_reg[16] [28]));
   NOR2_X1 i_4_0_590 (.A1(n_4_0_48), .A2(n_4_0_30), .ZN(\partial_reg[16] [29]));
   NOR2_X1 i_4_0_591 (.A1(n_4_0_48), .A2(n_4_0_31), .ZN(\partial_reg[16] [30]));
   NOR2_X1 i_4_0_592 (.A1(n_4_0_48), .A2(n_4_0_32), .ZN(\partial_reg[16] [31]));
   INV_X1 i_4_0_593 (.A(op2[17]), .ZN(n_4_0_49));
   NOR2_X1 i_4_0_594 (.A1(n_4_0_49), .A2(n_4_0_1), .ZN(\partial_reg[17] [0]));
   NOR2_X1 i_4_0_595 (.A1(n_4_0_49), .A2(n_4_0_2), .ZN(\partial_reg[17] [1]));
   NOR2_X1 i_4_0_596 (.A1(n_4_0_49), .A2(n_4_0_3), .ZN(\partial_reg[17] [2]));
   NOR2_X1 i_4_0_597 (.A1(n_4_0_49), .A2(n_4_0_4), .ZN(\partial_reg[17] [3]));
   NOR2_X1 i_4_0_598 (.A1(n_4_0_49), .A2(n_4_0_5), .ZN(\partial_reg[17] [4]));
   NOR2_X1 i_4_0_599 (.A1(n_4_0_49), .A2(n_4_0_6), .ZN(\partial_reg[17] [5]));
   NOR2_X1 i_4_0_600 (.A1(n_4_0_49), .A2(n_4_0_7), .ZN(\partial_reg[17] [6]));
   NOR2_X1 i_4_0_601 (.A1(n_4_0_49), .A2(n_4_0_8), .ZN(\partial_reg[17] [7]));
   NOR2_X1 i_4_0_602 (.A1(n_4_0_49), .A2(n_4_0_9), .ZN(\partial_reg[17] [8]));
   NOR2_X1 i_4_0_603 (.A1(n_4_0_49), .A2(n_4_0_10), .ZN(\partial_reg[17] [9]));
   NOR2_X1 i_4_0_604 (.A1(n_4_0_49), .A2(n_4_0_11), .ZN(\partial_reg[17] [10]));
   NOR2_X1 i_4_0_605 (.A1(n_4_0_49), .A2(n_4_0_12), .ZN(\partial_reg[17] [11]));
   NOR2_X1 i_4_0_606 (.A1(n_4_0_49), .A2(n_4_0_13), .ZN(\partial_reg[17] [12]));
   NOR2_X1 i_4_0_607 (.A1(n_4_0_49), .A2(n_4_0_14), .ZN(\partial_reg[17] [13]));
   NOR2_X1 i_4_0_608 (.A1(n_4_0_49), .A2(n_4_0_15), .ZN(\partial_reg[17] [14]));
   NOR2_X1 i_4_0_609 (.A1(n_4_0_49), .A2(n_4_0_16), .ZN(\partial_reg[17] [15]));
   NOR2_X1 i_4_0_610 (.A1(n_4_0_49), .A2(n_4_0_17), .ZN(\partial_reg[17] [16]));
   NOR2_X1 i_4_0_611 (.A1(n_4_0_49), .A2(n_4_0_18), .ZN(\partial_reg[17] [17]));
   NOR2_X1 i_4_0_612 (.A1(n_4_0_49), .A2(n_4_0_19), .ZN(\partial_reg[17] [18]));
   NOR2_X1 i_4_0_613 (.A1(n_4_0_49), .A2(n_4_0_20), .ZN(\partial_reg[17] [19]));
   NOR2_X1 i_4_0_614 (.A1(n_4_0_49), .A2(n_4_0_21), .ZN(\partial_reg[17] [20]));
   NOR2_X1 i_4_0_615 (.A1(n_4_0_49), .A2(n_4_0_22), .ZN(\partial_reg[17] [21]));
   NOR2_X1 i_4_0_616 (.A1(n_4_0_49), .A2(n_4_0_23), .ZN(\partial_reg[17] [22]));
   NOR2_X1 i_4_0_617 (.A1(n_4_0_49), .A2(n_4_0_24), .ZN(\partial_reg[17] [23]));
   NOR2_X1 i_4_0_618 (.A1(n_4_0_49), .A2(n_4_0_25), .ZN(\partial_reg[17] [24]));
   NOR2_X1 i_4_0_619 (.A1(n_4_0_49), .A2(n_4_0_26), .ZN(\partial_reg[17] [25]));
   NOR2_X1 i_4_0_620 (.A1(n_4_0_49), .A2(n_4_0_27), .ZN(\partial_reg[17] [26]));
   NOR2_X1 i_4_0_621 (.A1(n_4_0_49), .A2(n_4_0_28), .ZN(\partial_reg[17] [27]));
   NOR2_X1 i_4_0_622 (.A1(n_4_0_49), .A2(n_4_0_29), .ZN(\partial_reg[17] [28]));
   NOR2_X1 i_4_0_623 (.A1(n_4_0_49), .A2(n_4_0_30), .ZN(\partial_reg[17] [29]));
   NOR2_X1 i_4_0_624 (.A1(n_4_0_49), .A2(n_4_0_31), .ZN(\partial_reg[17] [30]));
   NOR2_X1 i_4_0_625 (.A1(n_4_0_49), .A2(n_4_0_32), .ZN(\partial_reg[17] [31]));
   INV_X1 i_4_0_626 (.A(op2[18]), .ZN(n_4_0_50));
   NOR2_X1 i_4_0_627 (.A1(n_4_0_50), .A2(n_4_0_1), .ZN(\partial_reg[18] [0]));
   NOR2_X1 i_4_0_628 (.A1(n_4_0_50), .A2(n_4_0_2), .ZN(\partial_reg[18] [1]));
   NOR2_X1 i_4_0_629 (.A1(n_4_0_50), .A2(n_4_0_3), .ZN(\partial_reg[18] [2]));
   NOR2_X1 i_4_0_630 (.A1(n_4_0_50), .A2(n_4_0_4), .ZN(\partial_reg[18] [3]));
   NOR2_X1 i_4_0_631 (.A1(n_4_0_50), .A2(n_4_0_5), .ZN(\partial_reg[18] [4]));
   NOR2_X1 i_4_0_632 (.A1(n_4_0_50), .A2(n_4_0_6), .ZN(\partial_reg[18] [5]));
   NOR2_X1 i_4_0_633 (.A1(n_4_0_50), .A2(n_4_0_7), .ZN(\partial_reg[18] [6]));
   NOR2_X1 i_4_0_634 (.A1(n_4_0_50), .A2(n_4_0_8), .ZN(\partial_reg[18] [7]));
   NOR2_X1 i_4_0_635 (.A1(n_4_0_50), .A2(n_4_0_9), .ZN(\partial_reg[18] [8]));
   NOR2_X1 i_4_0_636 (.A1(n_4_0_50), .A2(n_4_0_10), .ZN(\partial_reg[18] [9]));
   NOR2_X1 i_4_0_637 (.A1(n_4_0_50), .A2(n_4_0_11), .ZN(\partial_reg[18] [10]));
   NOR2_X1 i_4_0_638 (.A1(n_4_0_50), .A2(n_4_0_12), .ZN(\partial_reg[18] [11]));
   NOR2_X1 i_4_0_639 (.A1(n_4_0_50), .A2(n_4_0_13), .ZN(\partial_reg[18] [12]));
   NOR2_X1 i_4_0_640 (.A1(n_4_0_50), .A2(n_4_0_14), .ZN(\partial_reg[18] [13]));
   NOR2_X1 i_4_0_641 (.A1(n_4_0_50), .A2(n_4_0_15), .ZN(\partial_reg[18] [14]));
   NOR2_X1 i_4_0_642 (.A1(n_4_0_50), .A2(n_4_0_16), .ZN(\partial_reg[18] [15]));
   NOR2_X1 i_4_0_643 (.A1(n_4_0_50), .A2(n_4_0_17), .ZN(\partial_reg[18] [16]));
   NOR2_X1 i_4_0_644 (.A1(n_4_0_50), .A2(n_4_0_18), .ZN(\partial_reg[18] [17]));
   NOR2_X1 i_4_0_645 (.A1(n_4_0_50), .A2(n_4_0_19), .ZN(\partial_reg[18] [18]));
   NOR2_X1 i_4_0_646 (.A1(n_4_0_50), .A2(n_4_0_20), .ZN(\partial_reg[18] [19]));
   NOR2_X1 i_4_0_647 (.A1(n_4_0_50), .A2(n_4_0_21), .ZN(\partial_reg[18] [20]));
   NOR2_X1 i_4_0_648 (.A1(n_4_0_50), .A2(n_4_0_22), .ZN(\partial_reg[18] [21]));
   NOR2_X1 i_4_0_649 (.A1(n_4_0_50), .A2(n_4_0_23), .ZN(\partial_reg[18] [22]));
   NOR2_X1 i_4_0_650 (.A1(n_4_0_50), .A2(n_4_0_24), .ZN(\partial_reg[18] [23]));
   NOR2_X1 i_4_0_651 (.A1(n_4_0_50), .A2(n_4_0_25), .ZN(\partial_reg[18] [24]));
   NOR2_X1 i_4_0_652 (.A1(n_4_0_50), .A2(n_4_0_26), .ZN(\partial_reg[18] [25]));
   NOR2_X1 i_4_0_653 (.A1(n_4_0_50), .A2(n_4_0_27), .ZN(\partial_reg[18] [26]));
   NOR2_X1 i_4_0_654 (.A1(n_4_0_50), .A2(n_4_0_28), .ZN(\partial_reg[18] [27]));
   NOR2_X1 i_4_0_655 (.A1(n_4_0_50), .A2(n_4_0_29), .ZN(\partial_reg[18] [28]));
   NOR2_X1 i_4_0_656 (.A1(n_4_0_50), .A2(n_4_0_30), .ZN(\partial_reg[18] [29]));
   NOR2_X1 i_4_0_657 (.A1(n_4_0_50), .A2(n_4_0_31), .ZN(\partial_reg[18] [30]));
   NOR2_X1 i_4_0_658 (.A1(n_4_0_50), .A2(n_4_0_32), .ZN(\partial_reg[18] [31]));
   INV_X1 i_4_0_659 (.A(op2[19]), .ZN(n_4_0_51));
   NOR2_X1 i_4_0_660 (.A1(n_4_0_51), .A2(n_4_0_1), .ZN(\partial_reg[19] [0]));
   NOR2_X1 i_4_0_661 (.A1(n_4_0_51), .A2(n_4_0_2), .ZN(\partial_reg[19] [1]));
   NOR2_X1 i_4_0_662 (.A1(n_4_0_51), .A2(n_4_0_3), .ZN(\partial_reg[19] [2]));
   NOR2_X1 i_4_0_663 (.A1(n_4_0_51), .A2(n_4_0_4), .ZN(\partial_reg[19] [3]));
   NOR2_X1 i_4_0_664 (.A1(n_4_0_51), .A2(n_4_0_5), .ZN(\partial_reg[19] [4]));
   NOR2_X1 i_4_0_665 (.A1(n_4_0_51), .A2(n_4_0_6), .ZN(\partial_reg[19] [5]));
   NOR2_X1 i_4_0_666 (.A1(n_4_0_51), .A2(n_4_0_7), .ZN(\partial_reg[19] [6]));
   NOR2_X1 i_4_0_667 (.A1(n_4_0_51), .A2(n_4_0_8), .ZN(\partial_reg[19] [7]));
   NOR2_X1 i_4_0_668 (.A1(n_4_0_51), .A2(n_4_0_9), .ZN(\partial_reg[19] [8]));
   NOR2_X1 i_4_0_669 (.A1(n_4_0_51), .A2(n_4_0_10), .ZN(\partial_reg[19] [9]));
   NOR2_X1 i_4_0_670 (.A1(n_4_0_51), .A2(n_4_0_11), .ZN(\partial_reg[19] [10]));
   NOR2_X1 i_4_0_671 (.A1(n_4_0_51), .A2(n_4_0_12), .ZN(\partial_reg[19] [11]));
   NOR2_X1 i_4_0_672 (.A1(n_4_0_51), .A2(n_4_0_13), .ZN(\partial_reg[19] [12]));
   NOR2_X1 i_4_0_673 (.A1(n_4_0_51), .A2(n_4_0_14), .ZN(\partial_reg[19] [13]));
   NOR2_X1 i_4_0_674 (.A1(n_4_0_51), .A2(n_4_0_15), .ZN(\partial_reg[19] [14]));
   NOR2_X1 i_4_0_675 (.A1(n_4_0_51), .A2(n_4_0_16), .ZN(\partial_reg[19] [15]));
   NOR2_X1 i_4_0_676 (.A1(n_4_0_51), .A2(n_4_0_17), .ZN(\partial_reg[19] [16]));
   NOR2_X1 i_4_0_677 (.A1(n_4_0_51), .A2(n_4_0_18), .ZN(\partial_reg[19] [17]));
   NOR2_X1 i_4_0_678 (.A1(n_4_0_51), .A2(n_4_0_19), .ZN(\partial_reg[19] [18]));
   NOR2_X1 i_4_0_679 (.A1(n_4_0_51), .A2(n_4_0_20), .ZN(\partial_reg[19] [19]));
   NOR2_X1 i_4_0_680 (.A1(n_4_0_51), .A2(n_4_0_21), .ZN(\partial_reg[19] [20]));
   NOR2_X1 i_4_0_681 (.A1(n_4_0_51), .A2(n_4_0_22), .ZN(\partial_reg[19] [21]));
   NOR2_X1 i_4_0_682 (.A1(n_4_0_51), .A2(n_4_0_23), .ZN(\partial_reg[19] [22]));
   NOR2_X1 i_4_0_683 (.A1(n_4_0_51), .A2(n_4_0_24), .ZN(\partial_reg[19] [23]));
   NOR2_X1 i_4_0_684 (.A1(n_4_0_51), .A2(n_4_0_25), .ZN(\partial_reg[19] [24]));
   NOR2_X1 i_4_0_685 (.A1(n_4_0_51), .A2(n_4_0_26), .ZN(\partial_reg[19] [25]));
   NOR2_X1 i_4_0_686 (.A1(n_4_0_51), .A2(n_4_0_27), .ZN(\partial_reg[19] [26]));
   NOR2_X1 i_4_0_687 (.A1(n_4_0_51), .A2(n_4_0_28), .ZN(\partial_reg[19] [27]));
   NOR2_X1 i_4_0_688 (.A1(n_4_0_51), .A2(n_4_0_29), .ZN(\partial_reg[19] [28]));
   NOR2_X1 i_4_0_689 (.A1(n_4_0_51), .A2(n_4_0_30), .ZN(\partial_reg[19] [29]));
   NOR2_X1 i_4_0_690 (.A1(n_4_0_51), .A2(n_4_0_31), .ZN(\partial_reg[19] [30]));
   NOR2_X1 i_4_0_691 (.A1(n_4_0_51), .A2(n_4_0_32), .ZN(\partial_reg[19] [31]));
   INV_X1 i_4_0_692 (.A(op2[20]), .ZN(n_4_0_52));
   NOR2_X1 i_4_0_693 (.A1(n_4_0_52), .A2(n_4_0_1), .ZN(\partial_reg[20] [0]));
   NOR2_X1 i_4_0_694 (.A1(n_4_0_52), .A2(n_4_0_2), .ZN(\partial_reg[20] [1]));
   NOR2_X1 i_4_0_695 (.A1(n_4_0_52), .A2(n_4_0_3), .ZN(\partial_reg[20] [2]));
   NOR2_X1 i_4_0_696 (.A1(n_4_0_52), .A2(n_4_0_4), .ZN(\partial_reg[20] [3]));
   NOR2_X1 i_4_0_697 (.A1(n_4_0_52), .A2(n_4_0_5), .ZN(\partial_reg[20] [4]));
   NOR2_X1 i_4_0_698 (.A1(n_4_0_52), .A2(n_4_0_6), .ZN(\partial_reg[20] [5]));
   NOR2_X1 i_4_0_699 (.A1(n_4_0_52), .A2(n_4_0_7), .ZN(\partial_reg[20] [6]));
   NOR2_X1 i_4_0_700 (.A1(n_4_0_52), .A2(n_4_0_8), .ZN(\partial_reg[20] [7]));
   NOR2_X1 i_4_0_701 (.A1(n_4_0_52), .A2(n_4_0_9), .ZN(\partial_reg[20] [8]));
   NOR2_X1 i_4_0_702 (.A1(n_4_0_52), .A2(n_4_0_10), .ZN(\partial_reg[20] [9]));
   NOR2_X1 i_4_0_703 (.A1(n_4_0_52), .A2(n_4_0_11), .ZN(\partial_reg[20] [10]));
   NOR2_X1 i_4_0_704 (.A1(n_4_0_52), .A2(n_4_0_12), .ZN(\partial_reg[20] [11]));
   NOR2_X1 i_4_0_705 (.A1(n_4_0_52), .A2(n_4_0_13), .ZN(\partial_reg[20] [12]));
   NOR2_X1 i_4_0_706 (.A1(n_4_0_52), .A2(n_4_0_14), .ZN(\partial_reg[20] [13]));
   NOR2_X1 i_4_0_707 (.A1(n_4_0_52), .A2(n_4_0_15), .ZN(\partial_reg[20] [14]));
   NOR2_X1 i_4_0_708 (.A1(n_4_0_52), .A2(n_4_0_16), .ZN(\partial_reg[20] [15]));
   NOR2_X1 i_4_0_709 (.A1(n_4_0_52), .A2(n_4_0_17), .ZN(\partial_reg[20] [16]));
   NOR2_X1 i_4_0_710 (.A1(n_4_0_52), .A2(n_4_0_18), .ZN(\partial_reg[20] [17]));
   NOR2_X1 i_4_0_711 (.A1(n_4_0_52), .A2(n_4_0_19), .ZN(\partial_reg[20] [18]));
   NOR2_X1 i_4_0_712 (.A1(n_4_0_52), .A2(n_4_0_20), .ZN(\partial_reg[20] [19]));
   NOR2_X1 i_4_0_713 (.A1(n_4_0_52), .A2(n_4_0_21), .ZN(\partial_reg[20] [20]));
   NOR2_X1 i_4_0_714 (.A1(n_4_0_52), .A2(n_4_0_22), .ZN(\partial_reg[20] [21]));
   NOR2_X1 i_4_0_715 (.A1(n_4_0_52), .A2(n_4_0_23), .ZN(\partial_reg[20] [22]));
   NOR2_X1 i_4_0_716 (.A1(n_4_0_52), .A2(n_4_0_24), .ZN(\partial_reg[20] [23]));
   NOR2_X1 i_4_0_717 (.A1(n_4_0_52), .A2(n_4_0_25), .ZN(\partial_reg[20] [24]));
   NOR2_X1 i_4_0_718 (.A1(n_4_0_52), .A2(n_4_0_26), .ZN(\partial_reg[20] [25]));
   NOR2_X1 i_4_0_719 (.A1(n_4_0_52), .A2(n_4_0_27), .ZN(\partial_reg[20] [26]));
   NOR2_X1 i_4_0_720 (.A1(n_4_0_52), .A2(n_4_0_28), .ZN(\partial_reg[20] [27]));
   NOR2_X1 i_4_0_721 (.A1(n_4_0_52), .A2(n_4_0_29), .ZN(\partial_reg[20] [28]));
   NOR2_X1 i_4_0_722 (.A1(n_4_0_52), .A2(n_4_0_30), .ZN(\partial_reg[20] [29]));
   NOR2_X1 i_4_0_723 (.A1(n_4_0_52), .A2(n_4_0_31), .ZN(\partial_reg[20] [30]));
   NOR2_X1 i_4_0_724 (.A1(n_4_0_52), .A2(n_4_0_32), .ZN(\partial_reg[20] [31]));
   INV_X1 i_4_0_725 (.A(op2[21]), .ZN(n_4_0_53));
   NOR2_X1 i_4_0_726 (.A1(n_4_0_53), .A2(n_4_0_1), .ZN(\partial_reg[21] [0]));
   NOR2_X1 i_4_0_727 (.A1(n_4_0_53), .A2(n_4_0_2), .ZN(\partial_reg[21] [1]));
   NOR2_X1 i_4_0_728 (.A1(n_4_0_53), .A2(n_4_0_3), .ZN(\partial_reg[21] [2]));
   NOR2_X1 i_4_0_729 (.A1(n_4_0_53), .A2(n_4_0_4), .ZN(\partial_reg[21] [3]));
   NOR2_X1 i_4_0_730 (.A1(n_4_0_53), .A2(n_4_0_5), .ZN(\partial_reg[21] [4]));
   NOR2_X1 i_4_0_731 (.A1(n_4_0_53), .A2(n_4_0_6), .ZN(\partial_reg[21] [5]));
   NOR2_X1 i_4_0_732 (.A1(n_4_0_53), .A2(n_4_0_7), .ZN(\partial_reg[21] [6]));
   NOR2_X1 i_4_0_733 (.A1(n_4_0_53), .A2(n_4_0_8), .ZN(\partial_reg[21] [7]));
   NOR2_X1 i_4_0_734 (.A1(n_4_0_53), .A2(n_4_0_9), .ZN(\partial_reg[21] [8]));
   NOR2_X1 i_4_0_735 (.A1(n_4_0_53), .A2(n_4_0_10), .ZN(\partial_reg[21] [9]));
   NOR2_X1 i_4_0_736 (.A1(n_4_0_53), .A2(n_4_0_11), .ZN(\partial_reg[21] [10]));
   NOR2_X1 i_4_0_737 (.A1(n_4_0_53), .A2(n_4_0_12), .ZN(\partial_reg[21] [11]));
   NOR2_X1 i_4_0_738 (.A1(n_4_0_53), .A2(n_4_0_13), .ZN(\partial_reg[21] [12]));
   NOR2_X1 i_4_0_739 (.A1(n_4_0_53), .A2(n_4_0_14), .ZN(\partial_reg[21] [13]));
   NOR2_X1 i_4_0_740 (.A1(n_4_0_53), .A2(n_4_0_15), .ZN(\partial_reg[21] [14]));
   NOR2_X1 i_4_0_741 (.A1(n_4_0_53), .A2(n_4_0_16), .ZN(\partial_reg[21] [15]));
   NOR2_X1 i_4_0_742 (.A1(n_4_0_53), .A2(n_4_0_17), .ZN(\partial_reg[21] [16]));
   NOR2_X1 i_4_0_743 (.A1(n_4_0_53), .A2(n_4_0_18), .ZN(\partial_reg[21] [17]));
   NOR2_X1 i_4_0_744 (.A1(n_4_0_53), .A2(n_4_0_19), .ZN(\partial_reg[21] [18]));
   NOR2_X1 i_4_0_745 (.A1(n_4_0_53), .A2(n_4_0_20), .ZN(\partial_reg[21] [19]));
   NOR2_X1 i_4_0_746 (.A1(n_4_0_53), .A2(n_4_0_21), .ZN(\partial_reg[21] [20]));
   NOR2_X1 i_4_0_747 (.A1(n_4_0_53), .A2(n_4_0_22), .ZN(\partial_reg[21] [21]));
   NOR2_X1 i_4_0_748 (.A1(n_4_0_53), .A2(n_4_0_23), .ZN(\partial_reg[21] [22]));
   NOR2_X1 i_4_0_749 (.A1(n_4_0_53), .A2(n_4_0_24), .ZN(\partial_reg[21] [23]));
   NOR2_X1 i_4_0_750 (.A1(n_4_0_53), .A2(n_4_0_25), .ZN(\partial_reg[21] [24]));
   NOR2_X1 i_4_0_751 (.A1(n_4_0_53), .A2(n_4_0_26), .ZN(\partial_reg[21] [25]));
   NOR2_X1 i_4_0_752 (.A1(n_4_0_53), .A2(n_4_0_27), .ZN(\partial_reg[21] [26]));
   NOR2_X1 i_4_0_753 (.A1(n_4_0_53), .A2(n_4_0_28), .ZN(\partial_reg[21] [27]));
   NOR2_X1 i_4_0_754 (.A1(n_4_0_53), .A2(n_4_0_29), .ZN(\partial_reg[21] [28]));
   NOR2_X1 i_4_0_755 (.A1(n_4_0_53), .A2(n_4_0_30), .ZN(\partial_reg[21] [29]));
   NOR2_X1 i_4_0_756 (.A1(n_4_0_53), .A2(n_4_0_31), .ZN(\partial_reg[21] [30]));
   NOR2_X1 i_4_0_757 (.A1(n_4_0_53), .A2(n_4_0_32), .ZN(\partial_reg[21] [31]));
   INV_X1 i_4_0_758 (.A(op2[22]), .ZN(n_4_0_54));
   NOR2_X1 i_4_0_759 (.A1(n_4_0_54), .A2(n_4_0_1), .ZN(\partial_reg[22] [0]));
   NOR2_X1 i_4_0_760 (.A1(n_4_0_54), .A2(n_4_0_2), .ZN(\partial_reg[22] [1]));
   NOR2_X1 i_4_0_761 (.A1(n_4_0_54), .A2(n_4_0_3), .ZN(\partial_reg[22] [2]));
   NOR2_X1 i_4_0_762 (.A1(n_4_0_54), .A2(n_4_0_4), .ZN(\partial_reg[22] [3]));
   NOR2_X1 i_4_0_763 (.A1(n_4_0_54), .A2(n_4_0_5), .ZN(\partial_reg[22] [4]));
   NOR2_X1 i_4_0_764 (.A1(n_4_0_54), .A2(n_4_0_6), .ZN(\partial_reg[22] [5]));
   NOR2_X1 i_4_0_765 (.A1(n_4_0_54), .A2(n_4_0_7), .ZN(\partial_reg[22] [6]));
   NOR2_X1 i_4_0_766 (.A1(n_4_0_54), .A2(n_4_0_8), .ZN(\partial_reg[22] [7]));
   NOR2_X1 i_4_0_767 (.A1(n_4_0_54), .A2(n_4_0_9), .ZN(\partial_reg[22] [8]));
   NOR2_X1 i_4_0_768 (.A1(n_4_0_54), .A2(n_4_0_10), .ZN(\partial_reg[22] [9]));
   NOR2_X1 i_4_0_769 (.A1(n_4_0_54), .A2(n_4_0_11), .ZN(\partial_reg[22] [10]));
   NOR2_X1 i_4_0_770 (.A1(n_4_0_54), .A2(n_4_0_12), .ZN(\partial_reg[22] [11]));
   NOR2_X1 i_4_0_771 (.A1(n_4_0_54), .A2(n_4_0_13), .ZN(\partial_reg[22] [12]));
   NOR2_X1 i_4_0_772 (.A1(n_4_0_54), .A2(n_4_0_14), .ZN(\partial_reg[22] [13]));
   NOR2_X1 i_4_0_773 (.A1(n_4_0_54), .A2(n_4_0_15), .ZN(\partial_reg[22] [14]));
   NOR2_X1 i_4_0_774 (.A1(n_4_0_54), .A2(n_4_0_16), .ZN(\partial_reg[22] [15]));
   NOR2_X1 i_4_0_775 (.A1(n_4_0_54), .A2(n_4_0_17), .ZN(\partial_reg[22] [16]));
   NOR2_X1 i_4_0_776 (.A1(n_4_0_54), .A2(n_4_0_18), .ZN(\partial_reg[22] [17]));
   NOR2_X1 i_4_0_777 (.A1(n_4_0_54), .A2(n_4_0_19), .ZN(\partial_reg[22] [18]));
   NOR2_X1 i_4_0_778 (.A1(n_4_0_54), .A2(n_4_0_20), .ZN(\partial_reg[22] [19]));
   NOR2_X1 i_4_0_779 (.A1(n_4_0_54), .A2(n_4_0_21), .ZN(\partial_reg[22] [20]));
   NOR2_X1 i_4_0_780 (.A1(n_4_0_54), .A2(n_4_0_22), .ZN(\partial_reg[22] [21]));
   NOR2_X1 i_4_0_781 (.A1(n_4_0_54), .A2(n_4_0_23), .ZN(\partial_reg[22] [22]));
   NOR2_X1 i_4_0_782 (.A1(n_4_0_54), .A2(n_4_0_24), .ZN(\partial_reg[22] [23]));
   NOR2_X1 i_4_0_783 (.A1(n_4_0_54), .A2(n_4_0_25), .ZN(\partial_reg[22] [24]));
   NOR2_X1 i_4_0_784 (.A1(n_4_0_54), .A2(n_4_0_26), .ZN(\partial_reg[22] [25]));
   NOR2_X1 i_4_0_785 (.A1(n_4_0_54), .A2(n_4_0_27), .ZN(\partial_reg[22] [26]));
   NOR2_X1 i_4_0_786 (.A1(n_4_0_54), .A2(n_4_0_28), .ZN(\partial_reg[22] [27]));
   NOR2_X1 i_4_0_787 (.A1(n_4_0_54), .A2(n_4_0_29), .ZN(\partial_reg[22] [28]));
   NOR2_X1 i_4_0_788 (.A1(n_4_0_54), .A2(n_4_0_30), .ZN(\partial_reg[22] [29]));
   NOR2_X1 i_4_0_789 (.A1(n_4_0_54), .A2(n_4_0_31), .ZN(\partial_reg[22] [30]));
   NOR2_X1 i_4_0_790 (.A1(n_4_0_54), .A2(n_4_0_32), .ZN(\partial_reg[22] [31]));
   INV_X1 i_4_0_791 (.A(op2[23]), .ZN(n_4_0_55));
   NOR2_X1 i_4_0_792 (.A1(n_4_0_55), .A2(n_4_0_1), .ZN(\partial_reg[23] [0]));
   NOR2_X1 i_4_0_793 (.A1(n_4_0_55), .A2(n_4_0_2), .ZN(\partial_reg[23] [1]));
   NOR2_X1 i_4_0_794 (.A1(n_4_0_55), .A2(n_4_0_3), .ZN(\partial_reg[23] [2]));
   NOR2_X1 i_4_0_795 (.A1(n_4_0_55), .A2(n_4_0_4), .ZN(\partial_reg[23] [3]));
   NOR2_X1 i_4_0_796 (.A1(n_4_0_55), .A2(n_4_0_5), .ZN(\partial_reg[23] [4]));
   NOR2_X1 i_4_0_797 (.A1(n_4_0_55), .A2(n_4_0_6), .ZN(\partial_reg[23] [5]));
   NOR2_X1 i_4_0_798 (.A1(n_4_0_55), .A2(n_4_0_7), .ZN(\partial_reg[23] [6]));
   NOR2_X1 i_4_0_799 (.A1(n_4_0_55), .A2(n_4_0_8), .ZN(\partial_reg[23] [7]));
   NOR2_X1 i_4_0_800 (.A1(n_4_0_55), .A2(n_4_0_9), .ZN(\partial_reg[23] [8]));
   NOR2_X1 i_4_0_801 (.A1(n_4_0_55), .A2(n_4_0_10), .ZN(\partial_reg[23] [9]));
   NOR2_X1 i_4_0_802 (.A1(n_4_0_55), .A2(n_4_0_11), .ZN(\partial_reg[23] [10]));
   NOR2_X1 i_4_0_803 (.A1(n_4_0_55), .A2(n_4_0_12), .ZN(\partial_reg[23] [11]));
   NOR2_X1 i_4_0_804 (.A1(n_4_0_55), .A2(n_4_0_13), .ZN(\partial_reg[23] [12]));
   NOR2_X1 i_4_0_805 (.A1(n_4_0_55), .A2(n_4_0_14), .ZN(\partial_reg[23] [13]));
   NOR2_X1 i_4_0_806 (.A1(n_4_0_55), .A2(n_4_0_15), .ZN(\partial_reg[23] [14]));
   NOR2_X1 i_4_0_807 (.A1(n_4_0_55), .A2(n_4_0_16), .ZN(\partial_reg[23] [15]));
   NOR2_X1 i_4_0_808 (.A1(n_4_0_55), .A2(n_4_0_17), .ZN(\partial_reg[23] [16]));
   NOR2_X1 i_4_0_809 (.A1(n_4_0_55), .A2(n_4_0_18), .ZN(\partial_reg[23] [17]));
   NOR2_X1 i_4_0_810 (.A1(n_4_0_55), .A2(n_4_0_19), .ZN(\partial_reg[23] [18]));
   NOR2_X1 i_4_0_811 (.A1(n_4_0_55), .A2(n_4_0_20), .ZN(\partial_reg[23] [19]));
   NOR2_X1 i_4_0_812 (.A1(n_4_0_55), .A2(n_4_0_21), .ZN(\partial_reg[23] [20]));
   NOR2_X1 i_4_0_813 (.A1(n_4_0_55), .A2(n_4_0_22), .ZN(\partial_reg[23] [21]));
   NOR2_X1 i_4_0_814 (.A1(n_4_0_55), .A2(n_4_0_23), .ZN(\partial_reg[23] [22]));
   NOR2_X1 i_4_0_815 (.A1(n_4_0_55), .A2(n_4_0_24), .ZN(\partial_reg[23] [23]));
   NOR2_X1 i_4_0_816 (.A1(n_4_0_55), .A2(n_4_0_25), .ZN(\partial_reg[23] [24]));
   NOR2_X1 i_4_0_817 (.A1(n_4_0_55), .A2(n_4_0_26), .ZN(\partial_reg[23] [25]));
   NOR2_X1 i_4_0_818 (.A1(n_4_0_55), .A2(n_4_0_27), .ZN(\partial_reg[23] [26]));
   NOR2_X1 i_4_0_819 (.A1(n_4_0_55), .A2(n_4_0_28), .ZN(\partial_reg[23] [27]));
   NOR2_X1 i_4_0_820 (.A1(n_4_0_55), .A2(n_4_0_29), .ZN(\partial_reg[23] [28]));
   NOR2_X1 i_4_0_821 (.A1(n_4_0_55), .A2(n_4_0_30), .ZN(\partial_reg[23] [29]));
   NOR2_X1 i_4_0_822 (.A1(n_4_0_55), .A2(n_4_0_31), .ZN(\partial_reg[23] [30]));
   NOR2_X1 i_4_0_823 (.A1(n_4_0_55), .A2(n_4_0_32), .ZN(\partial_reg[23] [31]));
   INV_X1 i_4_0_824 (.A(op2[24]), .ZN(n_4_0_56));
   NOR2_X1 i_4_0_825 (.A1(n_4_0_56), .A2(n_4_0_1), .ZN(\partial_reg[24] [0]));
   NOR2_X1 i_4_0_826 (.A1(n_4_0_56), .A2(n_4_0_2), .ZN(\partial_reg[24] [1]));
   NOR2_X1 i_4_0_827 (.A1(n_4_0_56), .A2(n_4_0_3), .ZN(\partial_reg[24] [2]));
   NOR2_X1 i_4_0_828 (.A1(n_4_0_56), .A2(n_4_0_4), .ZN(\partial_reg[24] [3]));
   NOR2_X1 i_4_0_829 (.A1(n_4_0_56), .A2(n_4_0_5), .ZN(\partial_reg[24] [4]));
   NOR2_X1 i_4_0_830 (.A1(n_4_0_56), .A2(n_4_0_6), .ZN(\partial_reg[24] [5]));
   NOR2_X1 i_4_0_831 (.A1(n_4_0_56), .A2(n_4_0_7), .ZN(\partial_reg[24] [6]));
   NOR2_X1 i_4_0_832 (.A1(n_4_0_56), .A2(n_4_0_8), .ZN(\partial_reg[24] [7]));
   NOR2_X1 i_4_0_833 (.A1(n_4_0_56), .A2(n_4_0_9), .ZN(\partial_reg[24] [8]));
   NOR2_X1 i_4_0_834 (.A1(n_4_0_56), .A2(n_4_0_10), .ZN(\partial_reg[24] [9]));
   NOR2_X1 i_4_0_835 (.A1(n_4_0_56), .A2(n_4_0_11), .ZN(\partial_reg[24] [10]));
   NOR2_X1 i_4_0_836 (.A1(n_4_0_56), .A2(n_4_0_12), .ZN(\partial_reg[24] [11]));
   NOR2_X1 i_4_0_837 (.A1(n_4_0_56), .A2(n_4_0_13), .ZN(\partial_reg[24] [12]));
   NOR2_X1 i_4_0_838 (.A1(n_4_0_56), .A2(n_4_0_14), .ZN(\partial_reg[24] [13]));
   NOR2_X1 i_4_0_839 (.A1(n_4_0_56), .A2(n_4_0_15), .ZN(\partial_reg[24] [14]));
   NOR2_X1 i_4_0_840 (.A1(n_4_0_56), .A2(n_4_0_16), .ZN(\partial_reg[24] [15]));
   NOR2_X1 i_4_0_841 (.A1(n_4_0_56), .A2(n_4_0_17), .ZN(\partial_reg[24] [16]));
   NOR2_X1 i_4_0_842 (.A1(n_4_0_56), .A2(n_4_0_18), .ZN(\partial_reg[24] [17]));
   NOR2_X1 i_4_0_843 (.A1(n_4_0_56), .A2(n_4_0_19), .ZN(\partial_reg[24] [18]));
   NOR2_X1 i_4_0_844 (.A1(n_4_0_56), .A2(n_4_0_20), .ZN(\partial_reg[24] [19]));
   NOR2_X1 i_4_0_845 (.A1(n_4_0_56), .A2(n_4_0_21), .ZN(\partial_reg[24] [20]));
   NOR2_X1 i_4_0_846 (.A1(n_4_0_56), .A2(n_4_0_22), .ZN(\partial_reg[24] [21]));
   NOR2_X1 i_4_0_847 (.A1(n_4_0_56), .A2(n_4_0_23), .ZN(\partial_reg[24] [22]));
   NOR2_X1 i_4_0_848 (.A1(n_4_0_56), .A2(n_4_0_24), .ZN(\partial_reg[24] [23]));
   NOR2_X1 i_4_0_849 (.A1(n_4_0_56), .A2(n_4_0_25), .ZN(\partial_reg[24] [24]));
   NOR2_X1 i_4_0_850 (.A1(n_4_0_56), .A2(n_4_0_26), .ZN(\partial_reg[24] [25]));
   NOR2_X1 i_4_0_851 (.A1(n_4_0_56), .A2(n_4_0_27), .ZN(\partial_reg[24] [26]));
   NOR2_X1 i_4_0_852 (.A1(n_4_0_56), .A2(n_4_0_28), .ZN(\partial_reg[24] [27]));
   NOR2_X1 i_4_0_853 (.A1(n_4_0_56), .A2(n_4_0_29), .ZN(\partial_reg[24] [28]));
   NOR2_X1 i_4_0_854 (.A1(n_4_0_56), .A2(n_4_0_30), .ZN(\partial_reg[24] [29]));
   NOR2_X1 i_4_0_855 (.A1(n_4_0_56), .A2(n_4_0_31), .ZN(\partial_reg[24] [30]));
   NOR2_X1 i_4_0_856 (.A1(n_4_0_56), .A2(n_4_0_32), .ZN(\partial_reg[24] [31]));
   INV_X1 i_4_0_857 (.A(op2[25]), .ZN(n_4_0_57));
   NOR2_X1 i_4_0_858 (.A1(n_4_0_57), .A2(n_4_0_1), .ZN(\partial_reg[25] [0]));
   NOR2_X1 i_4_0_859 (.A1(n_4_0_57), .A2(n_4_0_2), .ZN(\partial_reg[25] [1]));
   NOR2_X1 i_4_0_860 (.A1(n_4_0_57), .A2(n_4_0_3), .ZN(\partial_reg[25] [2]));
   NOR2_X1 i_4_0_861 (.A1(n_4_0_57), .A2(n_4_0_4), .ZN(\partial_reg[25] [3]));
   NOR2_X1 i_4_0_862 (.A1(n_4_0_57), .A2(n_4_0_5), .ZN(\partial_reg[25] [4]));
   NOR2_X1 i_4_0_863 (.A1(n_4_0_57), .A2(n_4_0_6), .ZN(\partial_reg[25] [5]));
   NOR2_X1 i_4_0_864 (.A1(n_4_0_57), .A2(n_4_0_7), .ZN(\partial_reg[25] [6]));
   NOR2_X1 i_4_0_865 (.A1(n_4_0_57), .A2(n_4_0_8), .ZN(\partial_reg[25] [7]));
   NOR2_X1 i_4_0_866 (.A1(n_4_0_57), .A2(n_4_0_9), .ZN(\partial_reg[25] [8]));
   NOR2_X1 i_4_0_867 (.A1(n_4_0_57), .A2(n_4_0_10), .ZN(\partial_reg[25] [9]));
   NOR2_X1 i_4_0_868 (.A1(n_4_0_57), .A2(n_4_0_11), .ZN(\partial_reg[25] [10]));
   NOR2_X1 i_4_0_869 (.A1(n_4_0_57), .A2(n_4_0_12), .ZN(\partial_reg[25] [11]));
   NOR2_X1 i_4_0_870 (.A1(n_4_0_57), .A2(n_4_0_13), .ZN(\partial_reg[25] [12]));
   NOR2_X1 i_4_0_871 (.A1(n_4_0_57), .A2(n_4_0_14), .ZN(\partial_reg[25] [13]));
   NOR2_X1 i_4_0_872 (.A1(n_4_0_57), .A2(n_4_0_15), .ZN(\partial_reg[25] [14]));
   NOR2_X1 i_4_0_873 (.A1(n_4_0_57), .A2(n_4_0_16), .ZN(\partial_reg[25] [15]));
   NOR2_X1 i_4_0_874 (.A1(n_4_0_57), .A2(n_4_0_17), .ZN(\partial_reg[25] [16]));
   NOR2_X1 i_4_0_875 (.A1(n_4_0_57), .A2(n_4_0_18), .ZN(\partial_reg[25] [17]));
   NOR2_X1 i_4_0_876 (.A1(n_4_0_57), .A2(n_4_0_19), .ZN(\partial_reg[25] [18]));
   NOR2_X1 i_4_0_877 (.A1(n_4_0_57), .A2(n_4_0_20), .ZN(\partial_reg[25] [19]));
   NOR2_X1 i_4_0_878 (.A1(n_4_0_57), .A2(n_4_0_21), .ZN(\partial_reg[25] [20]));
   NOR2_X1 i_4_0_879 (.A1(n_4_0_57), .A2(n_4_0_22), .ZN(\partial_reg[25] [21]));
   NOR2_X1 i_4_0_880 (.A1(n_4_0_57), .A2(n_4_0_23), .ZN(\partial_reg[25] [22]));
   NOR2_X1 i_4_0_881 (.A1(n_4_0_57), .A2(n_4_0_24), .ZN(\partial_reg[25] [23]));
   NOR2_X1 i_4_0_882 (.A1(n_4_0_57), .A2(n_4_0_25), .ZN(\partial_reg[25] [24]));
   NOR2_X1 i_4_0_883 (.A1(n_4_0_57), .A2(n_4_0_26), .ZN(\partial_reg[25] [25]));
   NOR2_X1 i_4_0_884 (.A1(n_4_0_57), .A2(n_4_0_27), .ZN(\partial_reg[25] [26]));
   NOR2_X1 i_4_0_885 (.A1(n_4_0_57), .A2(n_4_0_28), .ZN(\partial_reg[25] [27]));
   NOR2_X1 i_4_0_886 (.A1(n_4_0_57), .A2(n_4_0_29), .ZN(\partial_reg[25] [28]));
   NOR2_X1 i_4_0_887 (.A1(n_4_0_57), .A2(n_4_0_30), .ZN(\partial_reg[25] [29]));
   NOR2_X1 i_4_0_888 (.A1(n_4_0_57), .A2(n_4_0_31), .ZN(\partial_reg[25] [30]));
   NOR2_X1 i_4_0_889 (.A1(n_4_0_57), .A2(n_4_0_32), .ZN(\partial_reg[25] [31]));
   INV_X1 i_4_0_890 (.A(op2[26]), .ZN(n_4_0_58));
   NOR2_X1 i_4_0_891 (.A1(n_4_0_58), .A2(n_4_0_1), .ZN(\partial_reg[26] [0]));
   NOR2_X1 i_4_0_892 (.A1(n_4_0_58), .A2(n_4_0_2), .ZN(\partial_reg[26] [1]));
   NOR2_X1 i_4_0_893 (.A1(n_4_0_58), .A2(n_4_0_3), .ZN(\partial_reg[26] [2]));
   NOR2_X1 i_4_0_894 (.A1(n_4_0_58), .A2(n_4_0_4), .ZN(\partial_reg[26] [3]));
   NOR2_X1 i_4_0_895 (.A1(n_4_0_58), .A2(n_4_0_5), .ZN(\partial_reg[26] [4]));
   NOR2_X1 i_4_0_896 (.A1(n_4_0_58), .A2(n_4_0_6), .ZN(\partial_reg[26] [5]));
   NOR2_X1 i_4_0_897 (.A1(n_4_0_58), .A2(n_4_0_7), .ZN(\partial_reg[26] [6]));
   NOR2_X1 i_4_0_898 (.A1(n_4_0_58), .A2(n_4_0_8), .ZN(\partial_reg[26] [7]));
   NOR2_X1 i_4_0_899 (.A1(n_4_0_58), .A2(n_4_0_9), .ZN(\partial_reg[26] [8]));
   NOR2_X1 i_4_0_900 (.A1(n_4_0_58), .A2(n_4_0_10), .ZN(\partial_reg[26] [9]));
   NOR2_X1 i_4_0_901 (.A1(n_4_0_58), .A2(n_4_0_11), .ZN(\partial_reg[26] [10]));
   NOR2_X1 i_4_0_902 (.A1(n_4_0_58), .A2(n_4_0_12), .ZN(\partial_reg[26] [11]));
   NOR2_X1 i_4_0_903 (.A1(n_4_0_58), .A2(n_4_0_13), .ZN(\partial_reg[26] [12]));
   NOR2_X1 i_4_0_904 (.A1(n_4_0_58), .A2(n_4_0_14), .ZN(\partial_reg[26] [13]));
   NOR2_X1 i_4_0_905 (.A1(n_4_0_58), .A2(n_4_0_15), .ZN(\partial_reg[26] [14]));
   NOR2_X1 i_4_0_906 (.A1(n_4_0_58), .A2(n_4_0_16), .ZN(\partial_reg[26] [15]));
   NOR2_X1 i_4_0_907 (.A1(n_4_0_58), .A2(n_4_0_17), .ZN(\partial_reg[26] [16]));
   NOR2_X1 i_4_0_908 (.A1(n_4_0_58), .A2(n_4_0_18), .ZN(\partial_reg[26] [17]));
   NOR2_X1 i_4_0_909 (.A1(n_4_0_58), .A2(n_4_0_19), .ZN(\partial_reg[26] [18]));
   NOR2_X1 i_4_0_910 (.A1(n_4_0_58), .A2(n_4_0_20), .ZN(\partial_reg[26] [19]));
   NOR2_X1 i_4_0_911 (.A1(n_4_0_58), .A2(n_4_0_21), .ZN(\partial_reg[26] [20]));
   NOR2_X1 i_4_0_912 (.A1(n_4_0_58), .A2(n_4_0_22), .ZN(\partial_reg[26] [21]));
   NOR2_X1 i_4_0_913 (.A1(n_4_0_58), .A2(n_4_0_23), .ZN(\partial_reg[26] [22]));
   NOR2_X1 i_4_0_914 (.A1(n_4_0_58), .A2(n_4_0_24), .ZN(\partial_reg[26] [23]));
   NOR2_X1 i_4_0_915 (.A1(n_4_0_58), .A2(n_4_0_25), .ZN(\partial_reg[26] [24]));
   NOR2_X1 i_4_0_916 (.A1(n_4_0_58), .A2(n_4_0_26), .ZN(\partial_reg[26] [25]));
   NOR2_X1 i_4_0_917 (.A1(n_4_0_58), .A2(n_4_0_27), .ZN(\partial_reg[26] [26]));
   NOR2_X1 i_4_0_918 (.A1(n_4_0_58), .A2(n_4_0_28), .ZN(\partial_reg[26] [27]));
   NOR2_X1 i_4_0_919 (.A1(n_4_0_58), .A2(n_4_0_29), .ZN(\partial_reg[26] [28]));
   NOR2_X1 i_4_0_920 (.A1(n_4_0_58), .A2(n_4_0_30), .ZN(\partial_reg[26] [29]));
   NOR2_X1 i_4_0_921 (.A1(n_4_0_58), .A2(n_4_0_31), .ZN(\partial_reg[26] [30]));
   NOR2_X1 i_4_0_922 (.A1(n_4_0_58), .A2(n_4_0_32), .ZN(\partial_reg[26] [31]));
   INV_X1 i_4_0_923 (.A(op2[27]), .ZN(n_4_0_59));
   NOR2_X1 i_4_0_924 (.A1(n_4_0_59), .A2(n_4_0_1), .ZN(\partial_reg[27] [0]));
   NOR2_X1 i_4_0_925 (.A1(n_4_0_59), .A2(n_4_0_2), .ZN(\partial_reg[27] [1]));
   NOR2_X1 i_4_0_926 (.A1(n_4_0_59), .A2(n_4_0_3), .ZN(\partial_reg[27] [2]));
   NOR2_X1 i_4_0_927 (.A1(n_4_0_59), .A2(n_4_0_4), .ZN(\partial_reg[27] [3]));
   NOR2_X1 i_4_0_928 (.A1(n_4_0_59), .A2(n_4_0_5), .ZN(\partial_reg[27] [4]));
   NOR2_X1 i_4_0_929 (.A1(n_4_0_59), .A2(n_4_0_6), .ZN(\partial_reg[27] [5]));
   NOR2_X1 i_4_0_930 (.A1(n_4_0_59), .A2(n_4_0_7), .ZN(\partial_reg[27] [6]));
   NOR2_X1 i_4_0_931 (.A1(n_4_0_59), .A2(n_4_0_8), .ZN(\partial_reg[27] [7]));
   NOR2_X1 i_4_0_932 (.A1(n_4_0_59), .A2(n_4_0_9), .ZN(\partial_reg[27] [8]));
   NOR2_X1 i_4_0_933 (.A1(n_4_0_59), .A2(n_4_0_10), .ZN(\partial_reg[27] [9]));
   NOR2_X1 i_4_0_934 (.A1(n_4_0_59), .A2(n_4_0_11), .ZN(\partial_reg[27] [10]));
   NOR2_X1 i_4_0_935 (.A1(n_4_0_59), .A2(n_4_0_12), .ZN(\partial_reg[27] [11]));
   NOR2_X1 i_4_0_936 (.A1(n_4_0_59), .A2(n_4_0_13), .ZN(\partial_reg[27] [12]));
   NOR2_X1 i_4_0_937 (.A1(n_4_0_59), .A2(n_4_0_14), .ZN(\partial_reg[27] [13]));
   NOR2_X1 i_4_0_938 (.A1(n_4_0_59), .A2(n_4_0_15), .ZN(\partial_reg[27] [14]));
   NOR2_X1 i_4_0_939 (.A1(n_4_0_59), .A2(n_4_0_16), .ZN(\partial_reg[27] [15]));
   NOR2_X1 i_4_0_940 (.A1(n_4_0_59), .A2(n_4_0_17), .ZN(\partial_reg[27] [16]));
   NOR2_X1 i_4_0_941 (.A1(n_4_0_59), .A2(n_4_0_18), .ZN(\partial_reg[27] [17]));
   NOR2_X1 i_4_0_942 (.A1(n_4_0_59), .A2(n_4_0_19), .ZN(\partial_reg[27] [18]));
   NOR2_X1 i_4_0_943 (.A1(n_4_0_59), .A2(n_4_0_20), .ZN(\partial_reg[27] [19]));
   NOR2_X1 i_4_0_944 (.A1(n_4_0_59), .A2(n_4_0_21), .ZN(\partial_reg[27] [20]));
   NOR2_X1 i_4_0_945 (.A1(n_4_0_59), .A2(n_4_0_22), .ZN(\partial_reg[27] [21]));
   NOR2_X1 i_4_0_946 (.A1(n_4_0_59), .A2(n_4_0_23), .ZN(\partial_reg[27] [22]));
   NOR2_X1 i_4_0_947 (.A1(n_4_0_59), .A2(n_4_0_24), .ZN(\partial_reg[27] [23]));
   NOR2_X1 i_4_0_948 (.A1(n_4_0_59), .A2(n_4_0_25), .ZN(\partial_reg[27] [24]));
   NOR2_X1 i_4_0_949 (.A1(n_4_0_59), .A2(n_4_0_26), .ZN(\partial_reg[27] [25]));
   NOR2_X1 i_4_0_950 (.A1(n_4_0_59), .A2(n_4_0_27), .ZN(\partial_reg[27] [26]));
   NOR2_X1 i_4_0_951 (.A1(n_4_0_59), .A2(n_4_0_28), .ZN(\partial_reg[27] [27]));
   NOR2_X1 i_4_0_952 (.A1(n_4_0_59), .A2(n_4_0_29), .ZN(\partial_reg[27] [28]));
   NOR2_X1 i_4_0_953 (.A1(n_4_0_59), .A2(n_4_0_30), .ZN(\partial_reg[27] [29]));
   NOR2_X1 i_4_0_954 (.A1(n_4_0_59), .A2(n_4_0_31), .ZN(\partial_reg[27] [30]));
   NOR2_X1 i_4_0_955 (.A1(n_4_0_59), .A2(n_4_0_32), .ZN(\partial_reg[27] [31]));
   INV_X1 i_4_0_956 (.A(op2[28]), .ZN(n_4_0_60));
   NOR2_X1 i_4_0_957 (.A1(n_4_0_60), .A2(n_4_0_1), .ZN(\partial_reg[28] [0]));
   NOR2_X1 i_4_0_958 (.A1(n_4_0_60), .A2(n_4_0_2), .ZN(\partial_reg[28] [1]));
   NOR2_X1 i_4_0_959 (.A1(n_4_0_60), .A2(n_4_0_3), .ZN(\partial_reg[28] [2]));
   NOR2_X1 i_4_0_960 (.A1(n_4_0_60), .A2(n_4_0_4), .ZN(\partial_reg[28] [3]));
   NOR2_X1 i_4_0_961 (.A1(n_4_0_60), .A2(n_4_0_5), .ZN(\partial_reg[28] [4]));
   NOR2_X1 i_4_0_962 (.A1(n_4_0_60), .A2(n_4_0_6), .ZN(\partial_reg[28] [5]));
   NOR2_X1 i_4_0_963 (.A1(n_4_0_60), .A2(n_4_0_7), .ZN(\partial_reg[28] [6]));
   NOR2_X1 i_4_0_964 (.A1(n_4_0_60), .A2(n_4_0_8), .ZN(\partial_reg[28] [7]));
   NOR2_X1 i_4_0_965 (.A1(n_4_0_60), .A2(n_4_0_9), .ZN(\partial_reg[28] [8]));
   NOR2_X1 i_4_0_966 (.A1(n_4_0_60), .A2(n_4_0_10), .ZN(\partial_reg[28] [9]));
   NOR2_X1 i_4_0_967 (.A1(n_4_0_60), .A2(n_4_0_11), .ZN(\partial_reg[28] [10]));
   NOR2_X1 i_4_0_968 (.A1(n_4_0_60), .A2(n_4_0_12), .ZN(\partial_reg[28] [11]));
   NOR2_X1 i_4_0_969 (.A1(n_4_0_60), .A2(n_4_0_13), .ZN(\partial_reg[28] [12]));
   NOR2_X1 i_4_0_970 (.A1(n_4_0_60), .A2(n_4_0_14), .ZN(\partial_reg[28] [13]));
   NOR2_X1 i_4_0_971 (.A1(n_4_0_60), .A2(n_4_0_15), .ZN(\partial_reg[28] [14]));
   NOR2_X1 i_4_0_972 (.A1(n_4_0_60), .A2(n_4_0_16), .ZN(\partial_reg[28] [15]));
   NOR2_X1 i_4_0_973 (.A1(n_4_0_60), .A2(n_4_0_17), .ZN(\partial_reg[28] [16]));
   NOR2_X1 i_4_0_974 (.A1(n_4_0_60), .A2(n_4_0_18), .ZN(\partial_reg[28] [17]));
   NOR2_X1 i_4_0_975 (.A1(n_4_0_60), .A2(n_4_0_19), .ZN(\partial_reg[28] [18]));
   NOR2_X1 i_4_0_976 (.A1(n_4_0_60), .A2(n_4_0_20), .ZN(\partial_reg[28] [19]));
   NOR2_X1 i_4_0_977 (.A1(n_4_0_60), .A2(n_4_0_21), .ZN(\partial_reg[28] [20]));
   NOR2_X1 i_4_0_978 (.A1(n_4_0_60), .A2(n_4_0_22), .ZN(\partial_reg[28] [21]));
   NOR2_X1 i_4_0_979 (.A1(n_4_0_60), .A2(n_4_0_23), .ZN(\partial_reg[28] [22]));
   NOR2_X1 i_4_0_980 (.A1(n_4_0_60), .A2(n_4_0_24), .ZN(\partial_reg[28] [23]));
   NOR2_X1 i_4_0_981 (.A1(n_4_0_60), .A2(n_4_0_25), .ZN(\partial_reg[28] [24]));
   NOR2_X1 i_4_0_982 (.A1(n_4_0_60), .A2(n_4_0_26), .ZN(\partial_reg[28] [25]));
   NOR2_X1 i_4_0_983 (.A1(n_4_0_60), .A2(n_4_0_27), .ZN(\partial_reg[28] [26]));
   NOR2_X1 i_4_0_984 (.A1(n_4_0_60), .A2(n_4_0_28), .ZN(\partial_reg[28] [27]));
   NOR2_X1 i_4_0_985 (.A1(n_4_0_60), .A2(n_4_0_29), .ZN(\partial_reg[28] [28]));
   NOR2_X1 i_4_0_986 (.A1(n_4_0_60), .A2(n_4_0_30), .ZN(\partial_reg[28] [29]));
   NOR2_X1 i_4_0_987 (.A1(n_4_0_60), .A2(n_4_0_31), .ZN(\partial_reg[28] [30]));
   NOR2_X1 i_4_0_988 (.A1(n_4_0_60), .A2(n_4_0_32), .ZN(\partial_reg[28] [31]));
   INV_X1 i_4_0_989 (.A(op2[29]), .ZN(n_4_0_61));
   NOR2_X1 i_4_0_990 (.A1(n_4_0_61), .A2(n_4_0_1), .ZN(\partial_reg[29] [0]));
   NOR2_X1 i_4_0_991 (.A1(n_4_0_61), .A2(n_4_0_2), .ZN(\partial_reg[29] [1]));
   NOR2_X1 i_4_0_992 (.A1(n_4_0_61), .A2(n_4_0_3), .ZN(\partial_reg[29] [2]));
   NOR2_X1 i_4_0_993 (.A1(n_4_0_61), .A2(n_4_0_4), .ZN(\partial_reg[29] [3]));
   NOR2_X1 i_4_0_994 (.A1(n_4_0_61), .A2(n_4_0_5), .ZN(\partial_reg[29] [4]));
   NOR2_X1 i_4_0_995 (.A1(n_4_0_61), .A2(n_4_0_6), .ZN(\partial_reg[29] [5]));
   NOR2_X1 i_4_0_996 (.A1(n_4_0_61), .A2(n_4_0_7), .ZN(\partial_reg[29] [6]));
   NOR2_X1 i_4_0_997 (.A1(n_4_0_61), .A2(n_4_0_8), .ZN(\partial_reg[29] [7]));
   NOR2_X1 i_4_0_998 (.A1(n_4_0_61), .A2(n_4_0_9), .ZN(\partial_reg[29] [8]));
   NOR2_X1 i_4_0_999 (.A1(n_4_0_61), .A2(n_4_0_10), .ZN(\partial_reg[29] [9]));
   NOR2_X1 i_4_0_1000 (.A1(n_4_0_61), .A2(n_4_0_11), .ZN(\partial_reg[29] [10]));
   NOR2_X1 i_4_0_1001 (.A1(n_4_0_61), .A2(n_4_0_12), .ZN(\partial_reg[29] [11]));
   NOR2_X1 i_4_0_1002 (.A1(n_4_0_61), .A2(n_4_0_13), .ZN(\partial_reg[29] [12]));
   NOR2_X1 i_4_0_1003 (.A1(n_4_0_61), .A2(n_4_0_14), .ZN(\partial_reg[29] [13]));
   NOR2_X1 i_4_0_1004 (.A1(n_4_0_61), .A2(n_4_0_15), .ZN(\partial_reg[29] [14]));
   NOR2_X1 i_4_0_1005 (.A1(n_4_0_61), .A2(n_4_0_16), .ZN(\partial_reg[29] [15]));
   NOR2_X1 i_4_0_1006 (.A1(n_4_0_61), .A2(n_4_0_17), .ZN(\partial_reg[29] [16]));
   NOR2_X1 i_4_0_1007 (.A1(n_4_0_61), .A2(n_4_0_18), .ZN(\partial_reg[29] [17]));
   NOR2_X1 i_4_0_1008 (.A1(n_4_0_61), .A2(n_4_0_19), .ZN(\partial_reg[29] [18]));
   NOR2_X1 i_4_0_1009 (.A1(n_4_0_61), .A2(n_4_0_20), .ZN(\partial_reg[29] [19]));
   NOR2_X1 i_4_0_1010 (.A1(n_4_0_61), .A2(n_4_0_21), .ZN(\partial_reg[29] [20]));
   NOR2_X1 i_4_0_1011 (.A1(n_4_0_61), .A2(n_4_0_22), .ZN(\partial_reg[29] [21]));
   NOR2_X1 i_4_0_1012 (.A1(n_4_0_61), .A2(n_4_0_23), .ZN(\partial_reg[29] [22]));
   NOR2_X1 i_4_0_1013 (.A1(n_4_0_61), .A2(n_4_0_24), .ZN(\partial_reg[29] [23]));
   NOR2_X1 i_4_0_1014 (.A1(n_4_0_61), .A2(n_4_0_25), .ZN(\partial_reg[29] [24]));
   NOR2_X1 i_4_0_1015 (.A1(n_4_0_61), .A2(n_4_0_26), .ZN(\partial_reg[29] [25]));
   NOR2_X1 i_4_0_1016 (.A1(n_4_0_61), .A2(n_4_0_27), .ZN(\partial_reg[29] [26]));
   NOR2_X1 i_4_0_1017 (.A1(n_4_0_61), .A2(n_4_0_28), .ZN(\partial_reg[29] [27]));
   NOR2_X1 i_4_0_1018 (.A1(n_4_0_61), .A2(n_4_0_29), .ZN(\partial_reg[29] [28]));
   NOR2_X1 i_4_0_1019 (.A1(n_4_0_61), .A2(n_4_0_30), .ZN(\partial_reg[29] [29]));
   NOR2_X1 i_4_0_1020 (.A1(n_4_0_61), .A2(n_4_0_31), .ZN(\partial_reg[29] [30]));
   NOR2_X1 i_4_0_1021 (.A1(n_4_0_61), .A2(n_4_0_32), .ZN(\partial_reg[29] [31]));
   INV_X1 i_4_0_1022 (.A(op2[30]), .ZN(n_4_0_62));
   NOR2_X1 i_4_0_1023 (.A1(n_4_0_62), .A2(n_4_0_1), .ZN(\partial_reg[30] [0]));
   NOR2_X1 i_4_0_1024 (.A1(n_4_0_62), .A2(n_4_0_2), .ZN(\partial_reg[30] [1]));
   NOR2_X1 i_4_0_1025 (.A1(n_4_0_62), .A2(n_4_0_3), .ZN(\partial_reg[30] [2]));
   NOR2_X1 i_4_0_1026 (.A1(n_4_0_62), .A2(n_4_0_4), .ZN(\partial_reg[30] [3]));
   NOR2_X1 i_4_0_1027 (.A1(n_4_0_62), .A2(n_4_0_5), .ZN(\partial_reg[30] [4]));
   NOR2_X1 i_4_0_1028 (.A1(n_4_0_62), .A2(n_4_0_6), .ZN(\partial_reg[30] [5]));
   NOR2_X1 i_4_0_1029 (.A1(n_4_0_62), .A2(n_4_0_7), .ZN(\partial_reg[30] [6]));
   NOR2_X1 i_4_0_1030 (.A1(n_4_0_62), .A2(n_4_0_8), .ZN(\partial_reg[30] [7]));
   NOR2_X1 i_4_0_1031 (.A1(n_4_0_62), .A2(n_4_0_9), .ZN(\partial_reg[30] [8]));
   NOR2_X1 i_4_0_1032 (.A1(n_4_0_62), .A2(n_4_0_10), .ZN(\partial_reg[30] [9]));
   NOR2_X1 i_4_0_1033 (.A1(n_4_0_62), .A2(n_4_0_11), .ZN(\partial_reg[30] [10]));
   NOR2_X1 i_4_0_1034 (.A1(n_4_0_62), .A2(n_4_0_12), .ZN(\partial_reg[30] [11]));
   NOR2_X1 i_4_0_1035 (.A1(n_4_0_62), .A2(n_4_0_13), .ZN(\partial_reg[30] [12]));
   NOR2_X1 i_4_0_1036 (.A1(n_4_0_62), .A2(n_4_0_14), .ZN(\partial_reg[30] [13]));
   NOR2_X1 i_4_0_1037 (.A1(n_4_0_62), .A2(n_4_0_15), .ZN(\partial_reg[30] [14]));
   NOR2_X1 i_4_0_1038 (.A1(n_4_0_62), .A2(n_4_0_16), .ZN(\partial_reg[30] [15]));
   NOR2_X1 i_4_0_1039 (.A1(n_4_0_62), .A2(n_4_0_17), .ZN(\partial_reg[30] [16]));
   NOR2_X1 i_4_0_1040 (.A1(n_4_0_62), .A2(n_4_0_18), .ZN(\partial_reg[30] [17]));
   NOR2_X1 i_4_0_1041 (.A1(n_4_0_62), .A2(n_4_0_19), .ZN(\partial_reg[30] [18]));
   NOR2_X1 i_4_0_1042 (.A1(n_4_0_62), .A2(n_4_0_20), .ZN(\partial_reg[30] [19]));
   NOR2_X1 i_4_0_1043 (.A1(n_4_0_62), .A2(n_4_0_21), .ZN(\partial_reg[30] [20]));
   NOR2_X1 i_4_0_1044 (.A1(n_4_0_62), .A2(n_4_0_22), .ZN(\partial_reg[30] [21]));
   NOR2_X1 i_4_0_1045 (.A1(n_4_0_62), .A2(n_4_0_23), .ZN(\partial_reg[30] [22]));
   NOR2_X1 i_4_0_1046 (.A1(n_4_0_62), .A2(n_4_0_24), .ZN(\partial_reg[30] [23]));
   NOR2_X1 i_4_0_1047 (.A1(n_4_0_62), .A2(n_4_0_25), .ZN(\partial_reg[30] [24]));
   NOR2_X1 i_4_0_1048 (.A1(n_4_0_62), .A2(n_4_0_26), .ZN(\partial_reg[30] [25]));
   NOR2_X1 i_4_0_1049 (.A1(n_4_0_62), .A2(n_4_0_27), .ZN(\partial_reg[30] [26]));
   NOR2_X1 i_4_0_1050 (.A1(n_4_0_62), .A2(n_4_0_28), .ZN(\partial_reg[30] [27]));
   NOR2_X1 i_4_0_1051 (.A1(n_4_0_62), .A2(n_4_0_29), .ZN(\partial_reg[30] [28]));
   NOR2_X1 i_4_0_1052 (.A1(n_4_0_62), .A2(n_4_0_30), .ZN(\partial_reg[30] [29]));
   NOR2_X1 i_4_0_1053 (.A1(n_4_0_62), .A2(n_4_0_31), .ZN(\partial_reg[30] [30]));
   NOR2_X1 i_4_0_1054 (.A1(n_4_0_62), .A2(n_4_0_32), .ZN(\partial_reg[30] [31]));
   INV_X1 i_4_0_1055 (.A(op2[31]), .ZN(n_4_0_63));
   NOR2_X1 i_4_0_1056 (.A1(n_4_0_1), .A2(n_4_0_63), .ZN(\partial_reg[31] [0]));
   NOR2_X1 i_4_0_1057 (.A1(n_4_0_2), .A2(n_4_0_63), .ZN(\partial_reg[31] [1]));
   NOR2_X1 i_4_0_1058 (.A1(n_4_0_3), .A2(n_4_0_63), .ZN(\partial_reg[31] [2]));
   NOR2_X1 i_4_0_1059 (.A1(n_4_0_4), .A2(n_4_0_63), .ZN(\partial_reg[31] [3]));
   NOR2_X1 i_4_0_1060 (.A1(n_4_0_5), .A2(n_4_0_63), .ZN(\partial_reg[31] [4]));
   NOR2_X1 i_4_0_1061 (.A1(n_4_0_6), .A2(n_4_0_63), .ZN(\partial_reg[31] [5]));
   NOR2_X1 i_4_0_1062 (.A1(n_4_0_7), .A2(n_4_0_63), .ZN(\partial_reg[31] [6]));
   NOR2_X1 i_4_0_1063 (.A1(n_4_0_8), .A2(n_4_0_63), .ZN(\partial_reg[31] [7]));
   NOR2_X1 i_4_0_1064 (.A1(n_4_0_9), .A2(n_4_0_63), .ZN(\partial_reg[31] [8]));
   NOR2_X1 i_4_0_1065 (.A1(n_4_0_10), .A2(n_4_0_63), .ZN(\partial_reg[31] [9]));
   NOR2_X1 i_4_0_1066 (.A1(n_4_0_11), .A2(n_4_0_63), .ZN(\partial_reg[31] [10]));
   NOR2_X1 i_4_0_1067 (.A1(n_4_0_12), .A2(n_4_0_63), .ZN(\partial_reg[31] [11]));
   NOR2_X1 i_4_0_1068 (.A1(n_4_0_13), .A2(n_4_0_63), .ZN(\partial_reg[31] [12]));
   NOR2_X1 i_4_0_1069 (.A1(n_4_0_14), .A2(n_4_0_63), .ZN(\partial_reg[31] [13]));
   NOR2_X1 i_4_0_1070 (.A1(n_4_0_15), .A2(n_4_0_63), .ZN(\partial_reg[31] [14]));
   NOR2_X1 i_4_0_1071 (.A1(n_4_0_16), .A2(n_4_0_63), .ZN(\partial_reg[31] [15]));
   NOR2_X1 i_4_0_1072 (.A1(n_4_0_17), .A2(n_4_0_63), .ZN(\partial_reg[31] [16]));
   NOR2_X1 i_4_0_1073 (.A1(n_4_0_18), .A2(n_4_0_63), .ZN(\partial_reg[31] [17]));
   NOR2_X1 i_4_0_1074 (.A1(n_4_0_19), .A2(n_4_0_63), .ZN(\partial_reg[31] [18]));
   NOR2_X1 i_4_0_1075 (.A1(n_4_0_20), .A2(n_4_0_63), .ZN(\partial_reg[31] [19]));
   NOR2_X1 i_4_0_1076 (.A1(n_4_0_21), .A2(n_4_0_63), .ZN(\partial_reg[31] [20]));
   NOR2_X1 i_4_0_1077 (.A1(n_4_0_22), .A2(n_4_0_63), .ZN(\partial_reg[31] [21]));
   NOR2_X1 i_4_0_1078 (.A1(n_4_0_23), .A2(n_4_0_63), .ZN(\partial_reg[31] [22]));
   NOR2_X1 i_4_0_1079 (.A1(n_4_0_24), .A2(n_4_0_63), .ZN(\partial_reg[31] [23]));
   NOR2_X1 i_4_0_1080 (.A1(n_4_0_25), .A2(n_4_0_63), .ZN(\partial_reg[31] [24]));
   NOR2_X1 i_4_0_1081 (.A1(n_4_0_26), .A2(n_4_0_63), .ZN(\partial_reg[31] [25]));
   NOR2_X1 i_4_0_1082 (.A1(n_4_0_27), .A2(n_4_0_63), .ZN(\partial_reg[31] [26]));
   NOR2_X1 i_4_0_1083 (.A1(n_4_0_28), .A2(n_4_0_63), .ZN(\partial_reg[31] [27]));
   NOR2_X1 i_4_0_1084 (.A1(n_4_0_29), .A2(n_4_0_63), .ZN(\partial_reg[31] [28]));
   NOR2_X1 i_4_0_1085 (.A1(n_4_0_30), .A2(n_4_0_63), .ZN(\partial_reg[31] [29]));
   NOR2_X1 i_4_0_1086 (.A1(n_4_0_31), .A2(n_4_0_63), .ZN(\partial_reg[31] [30]));
   NOR2_X1 i_4_0_1087 (.A1(n_4_0_32), .A2(n_4_0_63), .ZN(\partial_reg[31] [31]));
   INV_X1 i_4_0_0 (.A(op2[2]), .ZN(n_4_0_34));
   INV_X1 i_4_0_59 (.A(op2[1]), .ZN(n_4_0_33));
   INV_X1 i_4_0_61 (.A(op1[31]), .ZN(n_4_0_32));
   INV_X1 i_4_0_63 (.A(op1[30]), .ZN(n_4_0_31));
   INV_X1 i_4_0_64 (.A(op1[29]), .ZN(n_4_0_30));
   INV_X1 i_4_0_65 (.A(b[0]), .ZN(n_4_0_0));
   INV_X1 i_4_0_96 (.A(n_4_0_64), .ZN(\partial_reg[1] [30]));
   NAND2_X1 i_4_0_97 (.A1(op1[30]), .A2(op2[1]), .ZN(n_4_0_64));
   INV_X1 i_4_0_98 (.A(n_4_0_65), .ZN(\partial_reg[1] [31]));
   NAND2_X1 i_4_0_128 (.A1(op1[31]), .A2(op2[1]), .ZN(n_4_0_65));
   AND2_X1 i_4_0_129 (.A1(op1[31]), .A2(b[0]), .ZN(\partial_reg[0] [31]));
   AND2_X1 i_4_0_1088 (.A1(op1[29]), .A2(op2[2]), .ZN(\partial_reg[2] [29]));
   AND2_X1 i_4_0_1089 (.A1(op1[30]), .A2(op2[2]), .ZN(\partial_reg[2] [30]));
   PartialAdder p1 (.a({uc_87, \partial_reg[0] [31], \partial_reg[0] [30], 
      \partial_reg[0] [29], \partial_reg[0] [28], \partial_reg[0] [27], 
      \partial_reg[0] [26], \partial_reg[0] [25], \partial_reg[0] [24], 
      \partial_reg[0] [23], \partial_reg[0] [22], \partial_reg[0] [21], 
      \partial_reg[0] [20], \partial_reg[0] [19], \partial_reg[0] [18], 
      \partial_reg[0] [17], \partial_reg[0] [16], \partial_reg[0] [15], 
      \partial_reg[0] [14], \partial_reg[0] [13], \partial_reg[0] [12], 
      \partial_reg[0] [11], \partial_reg[0] [10], \partial_reg[0] [9], 
      \partial_reg[0] [8], \partial_reg[0] [7], \partial_reg[0] [6], 
      \partial_reg[0] [5], \partial_reg[0] [4], \partial_reg[0] [3], 
      \partial_reg[0] [2], \partial_reg[0] [1], uc_88}), .b(\partial_reg[1] ), 
      .c({uc_89, \partial_reg[2] [30], \partial_reg[2] [29], 
      \partial_reg[2] [28], \partial_reg[2] [27], \partial_reg[2] [26], 
      \partial_reg[2] [25], \partial_reg[2] [24], \partial_reg[2] [23], 
      \partial_reg[2] [22], \partial_reg[2] [21], \partial_reg[2] [20], 
      \partial_reg[2] [19], \partial_reg[2] [18], \partial_reg[2] [17], 
      \partial_reg[2] [16], \partial_reg[2] [15], \partial_reg[2] [14], 
      \partial_reg[2] [13], \partial_reg[2] [12], \partial_reg[2] [11], 
      \partial_reg[2] [10], \partial_reg[2] [9], \partial_reg[2] [8], 
      \partial_reg[2] [7], \partial_reg[2] [6], \partial_reg[2] [5], 
      \partial_reg[2] [4], \partial_reg[2] [3], \partial_reg[2] [2], 
      \partial_reg[2] [1], \partial_reg[2] [0]}), .s1({uc_90, \s1[0] [31], 
      \s1[0] [30], \s1[0] [29], \s1[0] [28], \s1[0] [27], \s1[0] [26], 
      \s1[0] [25], \s1[0] [24], \s1[0] [23], \s1[0] [22], \s1[0] [21], 
      \s1[0] [20], \s1[0] [19], \s1[0] [18], \s1[0] [17], \s1[0] [16], 
      \s1[0] [15], \s1[0] [14], \s1[0] [13], \s1[0] [12], \s1[0] [11], 
      \s1[0] [10], \s1[0] [9], \s1[0] [8], \s1[0] [7], \s1[0] [6], \s1[0] [5], 
      \s1[0] [4], \s1[0] [3], \s1[0] [2], \s1[0] [1], \s1[0] [0]}), .c1(\c1[0] ));
   datapath__0_4 i_0_2 (.p_0({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
      n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, 
      n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, 
      n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, uc_91}), .b(b));
   datapath__0_3 i_0_0 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_92}), .a(a));
   datapath__0_38 i_0_36 (.p_0({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, uc_93}), .sum1({n_28, n_60, 
      n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
      n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
      n_35, n_34, n_33, n_32, n_31, n_30, n_29, \s1[29] [0], n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
      n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, 
      \s1[0] [0], out[0]}));
   MUX2_X1 i_0_1_1 (.A(b[1]), .B(n_0_31), .S(b[31]), .Z(op2[1]));
   MUX2_X1 i_0_1_2 (.A(b[2]), .B(n_0_32), .S(b[31]), .Z(op2[2]));
   MUX2_X1 i_0_1_3 (.A(b[3]), .B(n_0_33), .S(b[31]), .Z(op2[3]));
   MUX2_X1 i_0_1_4 (.A(b[4]), .B(n_0_34), .S(b[31]), .Z(op2[4]));
   MUX2_X1 i_0_1_5 (.A(b[5]), .B(n_0_35), .S(b[31]), .Z(op2[5]));
   MUX2_X1 i_0_1_6 (.A(b[6]), .B(n_0_36), .S(b[31]), .Z(op2[6]));
   MUX2_X1 i_0_1_7 (.A(b[7]), .B(n_0_37), .S(b[31]), .Z(op2[7]));
   MUX2_X1 i_0_1_8 (.A(b[8]), .B(n_0_38), .S(b[31]), .Z(op2[8]));
   MUX2_X1 i_0_1_9 (.A(b[9]), .B(n_0_39), .S(b[31]), .Z(op2[9]));
   MUX2_X1 i_0_1_10 (.A(b[10]), .B(n_0_40), .S(b[31]), .Z(op2[10]));
   MUX2_X1 i_0_1_11 (.A(b[11]), .B(n_0_41), .S(b[31]), .Z(op2[11]));
   MUX2_X1 i_0_1_12 (.A(b[12]), .B(n_0_42), .S(b[31]), .Z(op2[12]));
   MUX2_X1 i_0_1_13 (.A(b[13]), .B(n_0_43), .S(b[31]), .Z(op2[13]));
   MUX2_X1 i_0_1_14 (.A(b[14]), .B(n_0_44), .S(b[31]), .Z(op2[14]));
   MUX2_X1 i_0_1_15 (.A(b[15]), .B(n_0_45), .S(b[31]), .Z(op2[15]));
   MUX2_X1 i_0_1_16 (.A(b[16]), .B(n_0_46), .S(b[31]), .Z(op2[16]));
   MUX2_X1 i_0_1_17 (.A(b[17]), .B(n_0_47), .S(b[31]), .Z(op2[17]));
   MUX2_X1 i_0_1_18 (.A(b[18]), .B(n_0_48), .S(b[31]), .Z(op2[18]));
   MUX2_X1 i_0_1_19 (.A(b[19]), .B(n_0_49), .S(b[31]), .Z(op2[19]));
   MUX2_X1 i_0_1_20 (.A(b[20]), .B(n_0_50), .S(b[31]), .Z(op2[20]));
   MUX2_X1 i_0_1_21 (.A(b[21]), .B(n_0_51), .S(b[31]), .Z(op2[21]));
   MUX2_X1 i_0_1_22 (.A(b[22]), .B(n_0_52), .S(b[31]), .Z(op2[22]));
   MUX2_X1 i_0_1_23 (.A(b[23]), .B(n_0_53), .S(b[31]), .Z(op2[23]));
   MUX2_X1 i_0_1_24 (.A(b[24]), .B(n_0_54), .S(b[31]), .Z(op2[24]));
   MUX2_X1 i_0_1_25 (.A(b[25]), .B(n_0_55), .S(b[31]), .Z(op2[25]));
   MUX2_X1 i_0_1_26 (.A(b[26]), .B(n_0_56), .S(b[31]), .Z(op2[26]));
   MUX2_X1 i_0_1_27 (.A(b[27]), .B(n_0_57), .S(b[31]), .Z(op2[27]));
   MUX2_X1 i_0_1_28 (.A(b[28]), .B(n_0_58), .S(b[31]), .Z(op2[28]));
   MUX2_X1 i_0_1_29 (.A(b[29]), .B(n_0_59), .S(b[31]), .Z(op2[29]));
   MUX2_X1 i_0_1_30 (.A(b[30]), .B(n_0_60), .S(b[31]), .Z(op2[30]));
   AND2_X1 i_0_1_31 (.A1(n_0_61), .A2(b[31]), .ZN(op2[31]));
   MUX2_X1 i_0_1_32 (.A(a[1]), .B(n_0_0), .S(a[31]), .Z(op1[1]));
   MUX2_X1 i_0_1_33 (.A(a[2]), .B(n_0_1), .S(a[31]), .Z(op1[2]));
   MUX2_X1 i_0_1_34 (.A(a[3]), .B(n_0_2), .S(a[31]), .Z(op1[3]));
   MUX2_X1 i_0_1_35 (.A(a[4]), .B(n_0_3), .S(a[31]), .Z(op1[4]));
   MUX2_X1 i_0_1_36 (.A(a[5]), .B(n_0_4), .S(a[31]), .Z(op1[5]));
   MUX2_X1 i_0_1_37 (.A(a[6]), .B(n_0_5), .S(a[31]), .Z(op1[6]));
   MUX2_X1 i_0_1_38 (.A(a[7]), .B(n_0_6), .S(a[31]), .Z(op1[7]));
   MUX2_X1 i_0_1_39 (.A(a[8]), .B(n_0_7), .S(a[31]), .Z(op1[8]));
   MUX2_X1 i_0_1_40 (.A(a[9]), .B(n_0_8), .S(a[31]), .Z(op1[9]));
   MUX2_X1 i_0_1_41 (.A(a[10]), .B(n_0_9), .S(a[31]), .Z(op1[10]));
   MUX2_X1 i_0_1_42 (.A(a[11]), .B(n_0_10), .S(a[31]), .Z(op1[11]));
   MUX2_X1 i_0_1_43 (.A(a[12]), .B(n_0_11), .S(a[31]), .Z(op1[12]));
   MUX2_X1 i_0_1_44 (.A(a[13]), .B(n_0_12), .S(a[31]), .Z(op1[13]));
   MUX2_X1 i_0_1_45 (.A(a[14]), .B(n_0_13), .S(a[31]), .Z(op1[14]));
   MUX2_X1 i_0_1_46 (.A(a[15]), .B(n_0_14), .S(a[31]), .Z(op1[15]));
   MUX2_X1 i_0_1_47 (.A(a[16]), .B(n_0_15), .S(a[31]), .Z(op1[16]));
   MUX2_X1 i_0_1_48 (.A(a[17]), .B(n_0_16), .S(a[31]), .Z(op1[17]));
   MUX2_X1 i_0_1_59 (.A(a[28]), .B(n_0_27), .S(a[31]), .Z(op1[28]));
   MUX2_X1 i_0_1_60 (.A(a[29]), .B(n_0_28), .S(a[31]), .Z(op1[29]));
   MUX2_X1 i_0_1_61 (.A(a[30]), .B(n_0_29), .S(a[31]), .Z(op1[30]));
   AND2_X1 i_0_1_62 (.A1(n_0_30), .A2(a[31]), .ZN(op1[31]));
   MUX2_X1 i_0_1_63 (.A(n_0_62), .B(\s1[0] [0]), .S(n_0_1_11), .Z(out[1]));
   MUX2_X1 i_0_1_64 (.A(n_0_63), .B(n_0), .S(n_0_1_11), .Z(out[2]));
   MUX2_X1 i_0_1_65 (.A(n_0_64), .B(n_1), .S(n_0_1_11), .Z(out[3]));
   MUX2_X1 i_0_1_66 (.A(n_0_65), .B(n_2), .S(n_0_1_11), .Z(out[4]));
   MUX2_X1 i_0_1_67 (.A(n_0_66), .B(n_3), .S(n_0_1_11), .Z(out[5]));
   MUX2_X1 i_0_1_68 (.A(n_0_67), .B(n_4), .S(n_0_1_11), .Z(out[6]));
   MUX2_X1 i_0_1_69 (.A(n_0_68), .B(n_5), .S(n_0_1_11), .Z(out[7]));
   MUX2_X1 i_0_1_70 (.A(n_0_69), .B(n_6), .S(n_0_1_11), .Z(out[8]));
   MUX2_X1 i_0_1_71 (.A(n_0_70), .B(n_7), .S(n_0_1_11), .Z(out[9]));
   MUX2_X1 i_0_1_72 (.A(n_0_71), .B(n_8), .S(n_0_1_11), .Z(out[10]));
   MUX2_X1 i_0_1_73 (.A(n_0_72), .B(n_9), .S(n_0_1_11), .Z(out[11]));
   MUX2_X1 i_0_1_74 (.A(n_0_73), .B(n_10), .S(n_0_1_11), .Z(out[12]));
   MUX2_X1 i_0_1_75 (.A(n_0_74), .B(n_11), .S(n_0_1_11), .Z(out[13]));
   MUX2_X1 i_0_1_76 (.A(n_0_75), .B(n_12), .S(n_0_1_11), .Z(out[14]));
   MUX2_X1 i_0_1_77 (.A(n_0_76), .B(n_13), .S(n_0_1_11), .Z(out[15]));
   MUX2_X1 i_0_1_78 (.A(n_0_77), .B(n_14), .S(n_0_1_11), .Z(out[16]));
   MUX2_X1 i_0_1_79 (.A(n_0_78), .B(n_15), .S(n_0_1_11), .Z(out[17]));
   MUX2_X1 i_0_1_80 (.A(n_0_79), .B(n_16), .S(n_0_1_11), .Z(out[18]));
   MUX2_X1 i_0_1_81 (.A(n_0_80), .B(n_17), .S(n_0_1_11), .Z(out[19]));
   MUX2_X1 i_0_1_82 (.A(n_0_81), .B(n_18), .S(n_0_1_11), .Z(out[20]));
   MUX2_X1 i_0_1_83 (.A(n_0_82), .B(n_19), .S(n_0_1_11), .Z(out[21]));
   MUX2_X1 i_0_1_84 (.A(n_0_83), .B(n_20), .S(n_0_1_11), .Z(out[22]));
   MUX2_X1 i_0_1_85 (.A(n_0_84), .B(n_21), .S(n_0_1_11), .Z(out[23]));
   MUX2_X1 i_0_1_86 (.A(n_0_85), .B(n_22), .S(n_0_1_11), .Z(out[24]));
   MUX2_X1 i_0_1_87 (.A(n_0_86), .B(n_23), .S(n_0_1_11), .Z(out[25]));
   MUX2_X1 i_0_1_88 (.A(n_0_87), .B(n_24), .S(n_0_1_11), .Z(out[26]));
   MUX2_X1 i_0_1_89 (.A(n_0_88), .B(n_25), .S(n_0_1_11), .Z(out[27]));
   MUX2_X1 i_0_1_90 (.A(n_0_89), .B(n_26), .S(n_0_1_11), .Z(out[28]));
   MUX2_X1 i_0_1_91 (.A(n_0_90), .B(n_27), .S(n_0_1_11), .Z(out[29]));
   MUX2_X1 i_0_1_92 (.A(n_0_91), .B(\s1[29] [0]), .S(n_0_1_11), .Z(out[30]));
   MUX2_X1 i_0_1_93 (.A(n_0_92), .B(n_29), .S(n_0_1_11), .Z(out[31]));
   MUX2_X1 i_0_1_94 (.A(n_0_93), .B(n_30), .S(n_0_1_11), .Z(out[32]));
   MUX2_X1 i_0_1_95 (.A(n_0_94), .B(n_31), .S(n_0_1_11), .Z(out[33]));
   MUX2_X1 i_0_1_96 (.A(n_0_95), .B(n_32), .S(n_0_1_11), .Z(out[34]));
   MUX2_X1 i_0_1_97 (.A(n_0_96), .B(n_33), .S(n_0_1_11), .Z(out[35]));
   MUX2_X1 i_0_1_98 (.A(n_0_97), .B(n_34), .S(n_0_1_11), .Z(out[36]));
   MUX2_X1 i_0_1_99 (.A(n_0_98), .B(n_35), .S(n_0_1_11), .Z(out[37]));
   MUX2_X1 i_0_1_100 (.A(n_0_99), .B(n_36), .S(n_0_1_11), .Z(out[38]));
   MUX2_X1 i_0_1_101 (.A(n_0_100), .B(n_37), .S(n_0_1_11), .Z(out[39]));
   MUX2_X1 i_0_1_102 (.A(n_0_101), .B(n_38), .S(n_0_1_11), .Z(out[40]));
   MUX2_X1 i_0_1_103 (.A(n_0_102), .B(n_39), .S(n_0_1_11), .Z(out[41]));
   MUX2_X1 i_0_1_104 (.A(n_0_103), .B(n_40), .S(n_0_1_11), .Z(out[42]));
   MUX2_X1 i_0_1_105 (.A(n_0_104), .B(n_41), .S(n_0_1_11), .Z(out[43]));
   MUX2_X1 i_0_1_106 (.A(n_0_105), .B(n_42), .S(n_0_1_11), .Z(out[44]));
   MUX2_X1 i_0_1_107 (.A(n_0_106), .B(n_43), .S(n_0_1_11), .Z(out[45]));
   MUX2_X1 i_0_1_108 (.A(n_0_107), .B(n_44), .S(n_0_1_11), .Z(out[46]));
   MUX2_X1 i_0_1_109 (.A(n_0_108), .B(n_45), .S(n_0_1_11), .Z(out[47]));
   MUX2_X1 i_0_1_110 (.A(n_0_109), .B(n_46), .S(n_0_1_11), .Z(out[48]));
   MUX2_X1 i_0_1_111 (.A(n_0_110), .B(n_47), .S(n_0_1_11), .Z(out[49]));
   MUX2_X1 i_0_1_112 (.A(n_0_111), .B(n_48), .S(n_0_1_11), .Z(out[50]));
   MUX2_X1 i_0_1_113 (.A(n_0_112), .B(n_49), .S(n_0_1_11), .Z(out[51]));
   MUX2_X1 i_0_1_114 (.A(n_0_113), .B(n_50), .S(n_0_1_11), .Z(out[52]));
   MUX2_X1 i_0_1_115 (.A(n_0_114), .B(n_51), .S(n_0_1_11), .Z(out[53]));
   MUX2_X1 i_0_1_116 (.A(n_0_115), .B(n_52), .S(n_0_1_11), .Z(out[54]));
   MUX2_X1 i_0_1_117 (.A(n_0_116), .B(n_53), .S(n_0_1_11), .Z(out[55]));
   MUX2_X1 i_0_1_118 (.A(n_0_117), .B(n_54), .S(n_0_1_11), .Z(out[56]));
   OAI21_X1 i_0_1_0 (.A(n_0_1_4), .B1(n_0_1_5), .B2(n_0_1_11), .ZN(out[57]));
   INV_X1 i_0_1_49 (.A(n_0_118), .ZN(n_0_1_5));
   MUX2_X1 i_0_1_124 (.A(n_0_119), .B(n_56), .S(n_0_1_11), .Z(out[58]));
   MUX2_X1 i_0_1_125 (.A(n_0_120), .B(n_57), .S(n_0_1_11), .Z(out[59]));
   MUX2_X1 i_0_1_126 (.A(n_0_121), .B(n_58), .S(n_0_1_11), .Z(out[60]));
   MUX2_X1 i_0_1_127 (.A(n_0_122), .B(n_59), .S(n_0_1_11), .Z(out[61]));
   OAI21_X1 i_0_1_50 (.A(n_0_1_6), .B1(n_0_1_7), .B2(n_0_1_11), .ZN(out[62]));
   NAND2_X1 i_0_1_51 (.A1(n_60), .A2(n_0_1_11), .ZN(n_0_1_6));
   INV_X1 i_0_1_52 (.A(n_0_123), .ZN(n_0_1_7));
   NAND2_X1 i_0_1_53 (.A1(n_0_1_9), .A2(n_0_1_8), .ZN(out[63]));
   NAND2_X1 i_0_1_54 (.A1(n_28), .A2(n_0_1_11), .ZN(n_0_1_8));
   NAND2_X1 i_0_1_55 (.A1(n_0_124), .A2(n_0_1_10), .ZN(n_0_1_9));
   INV_X1 i_0_1_56 (.A(n_0_1_11), .ZN(n_0_1_10));
   INV_X1 i_0_1_57 (.A(a[31]), .ZN(n_0_1_12));
   INV_X1 i_0_1_58 (.A(a[31]), .ZN(n_0_1_13));
   NAND2_X1 i_0_1_119 (.A1(n_0_1_14), .A2(n_0_1_15), .ZN(op1[18]));
   NAND2_X1 i_0_1_120 (.A1(n_0_1_0), .A2(a[18]), .ZN(n_0_1_14));
   NAND2_X1 i_0_1_121 (.A1(a[31]), .A2(n_0_17), .ZN(n_0_1_15));
   NAND2_X1 i_0_1_122 (.A1(n_0_1_16), .A2(n_0_1_17), .ZN(op1[19]));
   NAND2_X1 i_0_1_123 (.A1(n_0_1_0), .A2(a[19]), .ZN(n_0_1_16));
   NAND2_X1 i_0_1_128 (.A1(a[31]), .A2(n_0_18), .ZN(n_0_1_17));
   NAND2_X1 i_0_1_129 (.A1(n_0_1_19), .A2(n_0_1_18), .ZN(op1[20]));
   NAND2_X1 i_0_1_130 (.A1(a[20]), .A2(n_0_1_13), .ZN(n_0_1_18));
   NAND2_X1 i_0_1_131 (.A1(a[31]), .A2(n_0_19), .ZN(n_0_1_19));
   NAND2_X1 i_0_1_132 (.A1(n_0_1_20), .A2(n_0_1_21), .ZN(op1[21]));
   NAND2_X1 i_0_1_133 (.A1(n_0_1_0), .A2(a[21]), .ZN(n_0_1_20));
   NAND2_X1 i_0_1_134 (.A1(a[31]), .A2(n_0_20), .ZN(n_0_1_21));
   NAND2_X1 i_0_1_135 (.A1(n_0_1_22), .A2(n_0_1_23), .ZN(op1[23]));
   NAND2_X1 i_0_1_136 (.A1(n_0_1_0), .A2(a[23]), .ZN(n_0_1_22));
   NAND2_X1 i_0_1_137 (.A1(a[31]), .A2(n_0_22), .ZN(n_0_1_23));
   NAND2_X1 i_0_1_138 (.A1(n_0_1_25), .A2(n_0_1_24), .ZN(op1[24]));
   NAND2_X1 i_0_1_139 (.A1(a[24]), .A2(n_0_1_13), .ZN(n_0_1_24));
   NAND2_X1 i_0_1_140 (.A1(a[31]), .A2(n_0_23), .ZN(n_0_1_25));
   NAND2_X1 i_0_1_141 (.A1(n_0_1_26), .A2(n_0_1_27), .ZN(op1[25]));
   NAND2_X1 i_0_1_142 (.A1(n_0_1_0), .A2(a[25]), .ZN(n_0_1_26));
   NAND2_X1 i_0_1_143 (.A1(a[31]), .A2(n_0_24), .ZN(n_0_1_27));
   NAND2_X1 i_0_1_144 (.A1(n_0_1_28), .A2(n_0_1_29), .ZN(op1[26]));
   NAND2_X1 i_0_1_145 (.A1(n_0_1_0), .A2(a[26]), .ZN(n_0_1_28));
   NAND2_X1 i_0_1_146 (.A1(a[31]), .A2(n_0_25), .ZN(n_0_1_29));
   NAND2_X1 i_0_1_147 (.A1(n_0_1_30), .A2(n_0_1_1), .ZN(op1[27]));
   NAND2_X1 i_0_1_148 (.A1(n_0_1_0), .A2(a[27]), .ZN(n_0_1_30));
   INV_X1 i_0_1_149 (.A(a[31]), .ZN(n_0_1_0));
   NAND2_X1 i_0_1_150 (.A1(a[31]), .A2(n_0_26), .ZN(n_0_1_1));
   NAND2_X1 i_0_1_151 (.A1(n_0_1_2), .A2(n_0_1_3), .ZN(op1[22]));
   NAND2_X1 i_0_1_152 (.A1(n_0_21), .A2(a[31]), .ZN(n_0_1_2));
   NAND2_X1 i_0_1_153 (.A1(n_0_1_12), .A2(a[22]), .ZN(n_0_1_3));
   NAND2_X1 i_0_1_154 (.A1(n_55), .A2(n_0_1_11), .ZN(n_0_1_4));
   XNOR2_X1 i_0_1_155 (.A(b[31]), .B(a[31]), .ZN(n_0_1_11));
endmodule

module Register__5_0(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module Register(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module Register__parameterized0(in, clk, out);
   input [63:0]in;
   input clk;
   output [63:0]out;

   DFF_X1 \out_reg[63]  (.D(in[63]), .CK(clk), .Q(out[63]), .QN());
   DFF_X1 \out_reg[62]  (.D(in[62]), .CK(clk), .Q(out[62]), .QN());
   DFF_X1 \out_reg[61]  (.D(in[61]), .CK(clk), .Q(out[61]), .QN());
   DFF_X1 \out_reg[60]  (.D(in[60]), .CK(clk), .Q(out[60]), .QN());
   DFF_X1 \out_reg[59]  (.D(in[59]), .CK(clk), .Q(out[59]), .QN());
   DFF_X1 \out_reg[58]  (.D(in[58]), .CK(clk), .Q(out[58]), .QN());
   DFF_X1 \out_reg[57]  (.D(in[57]), .CK(clk), .Q(out[57]), .QN());
   DFF_X1 \out_reg[56]  (.D(in[56]), .CK(clk), .Q(out[56]), .QN());
   DFF_X1 \out_reg[55]  (.D(in[55]), .CK(clk), .Q(out[55]), .QN());
   DFF_X1 \out_reg[54]  (.D(in[54]), .CK(clk), .Q(out[54]), .QN());
   DFF_X1 \out_reg[53]  (.D(in[53]), .CK(clk), .Q(out[53]), .QN());
   DFF_X1 \out_reg[52]  (.D(in[52]), .CK(clk), .Q(out[52]), .QN());
   DFF_X1 \out_reg[51]  (.D(in[51]), .CK(clk), .Q(out[51]), .QN());
   DFF_X1 \out_reg[50]  (.D(in[50]), .CK(clk), .Q(out[50]), .QN());
   DFF_X1 \out_reg[49]  (.D(in[49]), .CK(clk), .Q(out[49]), .QN());
   DFF_X1 \out_reg[48]  (.D(in[48]), .CK(clk), .Q(out[48]), .QN());
   DFF_X1 \out_reg[47]  (.D(in[47]), .CK(clk), .Q(out[47]), .QN());
   DFF_X1 \out_reg[46]  (.D(in[46]), .CK(clk), .Q(out[46]), .QN());
   DFF_X1 \out_reg[45]  (.D(in[45]), .CK(clk), .Q(out[45]), .QN());
   DFF_X1 \out_reg[44]  (.D(in[44]), .CK(clk), .Q(out[44]), .QN());
   DFF_X1 \out_reg[43]  (.D(in[43]), .CK(clk), .Q(out[43]), .QN());
   DFF_X1 \out_reg[42]  (.D(in[42]), .CK(clk), .Q(out[42]), .QN());
   DFF_X1 \out_reg[41]  (.D(in[41]), .CK(clk), .Q(out[41]), .QN());
   DFF_X1 \out_reg[40]  (.D(in[40]), .CK(clk), .Q(out[40]), .QN());
   DFF_X1 \out_reg[39]  (.D(in[39]), .CK(clk), .Q(out[39]), .QN());
   DFF_X1 \out_reg[38]  (.D(in[38]), .CK(clk), .Q(out[38]), .QN());
   DFF_X1 \out_reg[37]  (.D(in[37]), .CK(clk), .Q(out[37]), .QN());
   DFF_X1 \out_reg[36]  (.D(in[36]), .CK(clk), .Q(out[36]), .QN());
   DFF_X1 \out_reg[35]  (.D(in[35]), .CK(clk), .Q(out[35]), .QN());
   DFF_X1 \out_reg[34]  (.D(in[34]), .CK(clk), .Q(out[34]), .QN());
   DFF_X1 \out_reg[33]  (.D(in[33]), .CK(clk), .Q(out[33]), .QN());
   DFF_X1 \out_reg[32]  (.D(in[32]), .CK(clk), .Q(out[32]), .QN());
   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module TreeMultiplier(a, b, clk, data);
   input [31:0]a;
   input [31:0]b;
   input clk;
   output [63:0]data;

   wire [63:0]out;
   wire [31:0]c;
   wire [31:0]d;

   TreeMultiplierCirc t1 (.a(c), .b(d), .out(out));
   Register__5_0 Register_inst1 (.in(a), .clk(clk), .out(c));
   Register Register_inst2 (.in(b), .clk(clk), .out(d));
   Register__parameterized0 Register_inst3 (.in(out), .clk(clk), .out(data));
endmodule
