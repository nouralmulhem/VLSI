/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 23 16:53:43 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 4261203052 */

module regFile__0_18(read_data, read_data2, write_en, write_data, write_data2, 
      clk);
   output [31:0]read_data;
   output [31:0]read_data2;
   input write_en;
   input [31:0]write_data;
   input [31:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[31]  (.D(write_data2[31]), .CK(n_0), .Q(read_data2[31]), 
      .QN());
   DFF_X1 \my_reg2_reg[30]  (.D(write_data2[30]), .CK(n_0), .Q(read_data2[30]), 
      .QN());
   DFF_X1 \my_reg2_reg[29]  (.D(write_data2[29]), .CK(n_0), .Q(read_data2[29]), 
      .QN());
   DFF_X1 \my_reg2_reg[28]  (.D(write_data2[28]), .CK(n_0), .Q(read_data2[28]), 
      .QN());
   DFF_X1 \my_reg2_reg[27]  (.D(write_data2[27]), .CK(n_0), .Q(read_data2[27]), 
      .QN());
   DFF_X1 \my_reg2_reg[26]  (.D(write_data2[26]), .CK(n_0), .Q(read_data2[26]), 
      .QN());
   DFF_X1 \my_reg2_reg[25]  (.D(write_data2[25]), .CK(n_0), .Q(read_data2[25]), 
      .QN());
   DFF_X1 \my_reg2_reg[24]  (.D(write_data2[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data2[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
   DFF_X1 \my_reg2_reg[22]  (.D(write_data2[22]), .CK(n_0), .Q(read_data2[22]), 
      .QN());
   DFF_X1 \my_reg2_reg[21]  (.D(write_data2[21]), .CK(n_0), .Q(read_data2[21]), 
      .QN());
   DFF_X1 \my_reg2_reg[20]  (.D(write_data2[20]), .CK(n_0), .Q(read_data2[20]), 
      .QN());
   DFF_X1 \my_reg2_reg[19]  (.D(write_data2[19]), .CK(n_0), .Q(read_data2[19]), 
      .QN());
   DFF_X1 \my_reg2_reg[18]  (.D(write_data2[18]), .CK(n_0), .Q(read_data2[18]), 
      .QN());
   DFF_X1 \my_reg2_reg[17]  (.D(write_data2[17]), .CK(n_0), .Q(read_data2[17]), 
      .QN());
   DFF_X1 \my_reg2_reg[16]  (.D(write_data2[16]), .CK(n_0), .Q(read_data2[16]), 
      .QN());
   DFF_X1 \my_reg2_reg[15]  (.D(write_data2[15]), .CK(n_0), .Q(read_data2[15]), 
      .QN());
   DFF_X1 \my_reg2_reg[14]  (.D(write_data2[14]), .CK(n_0), .Q(read_data2[14]), 
      .QN());
   DFF_X1 \my_reg2_reg[13]  (.D(write_data2[13]), .CK(n_0), .Q(read_data2[13]), 
      .QN());
   DFF_X1 \my_reg2_reg[12]  (.D(write_data2[12]), .CK(n_0), .Q(read_data2[12]), 
      .QN());
   DFF_X1 \my_reg2_reg[11]  (.D(write_data2[11]), .CK(n_0), .Q(read_data2[11]), 
      .QN());
   DFF_X1 \my_reg2_reg[10]  (.D(write_data2[10]), .CK(n_0), .Q(read_data2[10]), 
      .QN());
   DFF_X1 \my_reg2_reg[9]  (.D(write_data2[9]), .CK(n_0), .Q(read_data2[9]), 
      .QN());
   DFF_X1 \my_reg2_reg[8]  (.D(write_data2[8]), .CK(n_0), .Q(read_data2[8]), 
      .QN());
   DFF_X1 \my_reg2_reg[7]  (.D(write_data2[7]), .CK(n_0), .Q(read_data2[7]), 
      .QN());
   DFF_X1 \my_reg2_reg[6]  (.D(write_data2[6]), .CK(n_0), .Q(read_data2[6]), 
      .QN());
   DFF_X1 \my_reg2_reg[5]  (.D(write_data2[5]), .CK(n_0), .Q(read_data2[5]), 
      .QN());
   DFF_X1 \my_reg2_reg[4]  (.D(write_data2[4]), .CK(n_0), .Q(read_data2[4]), 
      .QN());
   DFF_X1 \my_reg2_reg[3]  (.D(write_data2[3]), .CK(n_0), .Q(read_data2[3]), 
      .QN());
   DFF_X1 \my_reg2_reg[2]  (.D(write_data2[2]), .CK(n_0), .Q(read_data2[2]), 
      .QN());
   DFF_X1 \my_reg2_reg[1]  (.D(write_data2[1]), .CK(n_0), .Q(read_data2[1]), 
      .QN());
   DFF_X1 \my_reg2_reg[0]  (.D(write_data2[0]), .CK(n_0), .Q(read_data2[0]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg2_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
endmodule

module fullAdder__0_399(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_393(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_390(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_387(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_384(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_381(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_378(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_375(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_372(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_369(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_366(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_363(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_360(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_357(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_354(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_351(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_348(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_345(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_342(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_339(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_336(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_333(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_330(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_327(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_324(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_321(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_318(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_315(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_312(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_309(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_306(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_303(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_300(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(y), .B(x), .Z(sum));
endmodule

module fullAdder__0_297(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_294(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_291(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_288(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_285(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_282(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_279(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_276(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_273(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_270(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_267(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_264(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_261(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_258(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_255(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_252(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_249(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_246(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_243(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_240(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_237(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_234(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_231(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_228(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_225(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_222(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_219(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_216(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_210(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(x), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(y), .ZN(sum));
endmodule

module carrySaveAdder__0_400(a, b, c, sum, cout);
   input [31:0]a;
   input [31:0]b;
   input [31:0]c;
   output [31:0]sum;
   output cout;

   wire [31:0]halfcarry;
   wire [31:0]halfcout;
   wire [31:0]halfsum;

   fullAdder__0_399 fulladder_f2 (.x(halfsum[1]), .y(halfcout[0]), .cin(), 
      .sum(sum[1]), .cout(halfcarry[0]));
   fullAdder__0_393 genblk1_0_fulladder_f1 (.x(a[0]), .y(b[0]), .cin(), .sum(
      sum[0]), .cout(halfcout[0]));
   fullAdder__0_390 genblk1_1_fulladder_f1 (.x(a[1]), .y(b[1]), .cin(), .sum(
      halfsum[1]), .cout(halfcout[1]));
   fullAdder__0_387 genblk1_2_fulladder_f1 (.x(a[2]), .y(b[2]), .cin(), .sum(
      halfsum[2]), .cout(halfcout[2]));
   fullAdder__0_384 genblk1_3_fulladder_f1 (.x(a[3]), .y(b[3]), .cin(), .sum(
      halfsum[3]), .cout(halfcout[3]));
   fullAdder__0_381 genblk1_4_fulladder_f1 (.x(a[4]), .y(b[4]), .cin(), .sum(
      halfsum[4]), .cout(halfcout[4]));
   fullAdder__0_378 genblk1_5_fulladder_f1 (.x(a[5]), .y(b[5]), .cin(), .sum(
      halfsum[5]), .cout(halfcout[5]));
   fullAdder__0_375 genblk1_6_fulladder_f1 (.x(a[6]), .y(b[6]), .cin(), .sum(
      halfsum[6]), .cout(halfcout[6]));
   fullAdder__0_372 genblk1_7_fulladder_f1 (.x(a[7]), .y(b[7]), .cin(), .sum(
      halfsum[7]), .cout(halfcout[7]));
   fullAdder__0_369 genblk1_8_fulladder_f1 (.x(a[8]), .y(b[8]), .cin(), .sum(
      halfsum[8]), .cout(halfcout[8]));
   fullAdder__0_366 genblk1_9_fulladder_f1 (.x(a[9]), .y(b[9]), .cin(), .sum(
      halfsum[9]), .cout(halfcout[9]));
   fullAdder__0_363 genblk1_10_fulladder_f1 (.x(a[10]), .y(b[10]), .cin(), 
      .sum(halfsum[10]), .cout(halfcout[10]));
   fullAdder__0_360 genblk1_11_fulladder_f1 (.x(a[11]), .y(b[11]), .cin(), 
      .sum(halfsum[11]), .cout(halfcout[11]));
   fullAdder__0_357 genblk1_12_fulladder_f1 (.x(a[12]), .y(b[12]), .cin(), 
      .sum(halfsum[12]), .cout(halfcout[12]));
   fullAdder__0_354 genblk1_13_fulladder_f1 (.x(a[13]), .y(b[13]), .cin(), 
      .sum(halfsum[13]), .cout(halfcout[13]));
   fullAdder__0_351 genblk1_14_fulladder_f1 (.x(a[14]), .y(b[14]), .cin(), 
      .sum(halfsum[14]), .cout(halfcout[14]));
   fullAdder__0_348 genblk1_15_fulladder_f1 (.x(a[15]), .y(b[15]), .cin(), 
      .sum(halfsum[15]), .cout(halfcout[15]));
   fullAdder__0_345 genblk1_16_fulladder_f1 (.x(a[16]), .y(b[16]), .cin(), 
      .sum(halfsum[16]), .cout(halfcout[16]));
   fullAdder__0_342 genblk1_17_fulladder_f1 (.x(a[17]), .y(b[17]), .cin(), 
      .sum(halfsum[17]), .cout(halfcout[17]));
   fullAdder__0_339 genblk1_18_fulladder_f1 (.x(a[18]), .y(b[18]), .cin(), 
      .sum(halfsum[18]), .cout(halfcout[18]));
   fullAdder__0_336 genblk1_19_fulladder_f1 (.x(a[19]), .y(b[19]), .cin(), 
      .sum(halfsum[19]), .cout(halfcout[19]));
   fullAdder__0_333 genblk1_20_fulladder_f1 (.x(a[20]), .y(b[20]), .cin(), 
      .sum(halfsum[20]), .cout(halfcout[20]));
   fullAdder__0_330 genblk1_21_fulladder_f1 (.x(a[21]), .y(b[21]), .cin(), 
      .sum(halfsum[21]), .cout(halfcout[21]));
   fullAdder__0_327 genblk1_22_fulladder_f1 (.x(a[22]), .y(b[22]), .cin(), 
      .sum(halfsum[22]), .cout(halfcout[22]));
   fullAdder__0_324 genblk1_23_fulladder_f1 (.x(a[23]), .y(b[23]), .cin(), 
      .sum(halfsum[23]), .cout(halfcout[23]));
   fullAdder__0_321 genblk1_24_fulladder_f1 (.x(a[24]), .y(b[24]), .cin(), 
      .sum(halfsum[24]), .cout(halfcout[24]));
   fullAdder__0_318 genblk1_25_fulladder_f1 (.x(a[25]), .y(b[25]), .cin(), 
      .sum(halfsum[25]), .cout(halfcout[25]));
   fullAdder__0_315 genblk1_26_fulladder_f1 (.x(a[26]), .y(b[26]), .cin(), 
      .sum(halfsum[26]), .cout(halfcout[26]));
   fullAdder__0_312 genblk1_27_fulladder_f1 (.x(a[27]), .y(b[27]), .cin(), 
      .sum(halfsum[27]), .cout(halfcout[27]));
   fullAdder__0_309 genblk1_28_fulladder_f1 (.x(a[28]), .y(b[28]), .cin(), 
      .sum(halfsum[28]), .cout(halfcout[28]));
   fullAdder__0_306 genblk1_29_fulladder_f1 (.x(a[29]), .y(b[29]), .cin(), 
      .sum(halfsum[29]), .cout(halfcout[29]));
   fullAdder__0_303 genblk1_30_fulladder_f1 (.x(a[30]), .y(b[30]), .cin(), 
      .sum(halfsum[30]), .cout(halfcout[30]));
   fullAdder__0_300 genblk1_31_fulladder_f1 (.x(a[31]), .y(b[31]), .cin(), 
      .sum(halfsum[31]), .cout());
   fullAdder__0_297 genblk2_1_f3 (.x(halfsum[2]), .y(halfcout[1]), .cin(
      halfcarry[0]), .sum(sum[2]), .cout(halfcarry[1]));
   fullAdder__0_294 genblk2_2_f3 (.x(halfsum[3]), .y(halfcout[2]), .cin(
      halfcarry[1]), .sum(sum[3]), .cout(halfcarry[2]));
   fullAdder__0_291 genblk2_3_f3 (.x(halfsum[4]), .y(halfcout[3]), .cin(
      halfcarry[2]), .sum(sum[4]), .cout(halfcarry[3]));
   fullAdder__0_288 genblk2_4_f3 (.x(halfsum[5]), .y(halfcout[4]), .cin(
      halfcarry[3]), .sum(sum[5]), .cout(halfcarry[4]));
   fullAdder__0_285 genblk2_5_f3 (.x(halfsum[6]), .y(halfcout[5]), .cin(
      halfcarry[4]), .sum(sum[6]), .cout(halfcarry[5]));
   fullAdder__0_282 genblk2_6_f3 (.x(halfsum[7]), .y(halfcout[6]), .cin(
      halfcarry[5]), .sum(sum[7]), .cout(halfcarry[6]));
   fullAdder__0_279 genblk2_7_f3 (.x(halfsum[8]), .y(halfcout[7]), .cin(
      halfcarry[6]), .sum(sum[8]), .cout(halfcarry[7]));
   fullAdder__0_276 genblk2_8_f3 (.x(halfsum[9]), .y(halfcout[8]), .cin(
      halfcarry[7]), .sum(sum[9]), .cout(halfcarry[8]));
   fullAdder__0_273 genblk2_9_f3 (.x(halfsum[10]), .y(halfcout[9]), .cin(
      halfcarry[8]), .sum(sum[10]), .cout(halfcarry[9]));
   fullAdder__0_270 genblk2_10_f3 (.x(halfsum[11]), .y(halfcout[10]), .cin(
      halfcarry[9]), .sum(sum[11]), .cout(halfcarry[10]));
   fullAdder__0_267 genblk2_11_f3 (.x(halfsum[12]), .y(halfcout[11]), .cin(
      halfcarry[10]), .sum(sum[12]), .cout(halfcarry[11]));
   fullAdder__0_264 genblk2_12_f3 (.x(halfsum[13]), .y(halfcout[12]), .cin(
      halfcarry[11]), .sum(sum[13]), .cout(halfcarry[12]));
   fullAdder__0_261 genblk2_13_f3 (.x(halfsum[14]), .y(halfcout[13]), .cin(
      halfcarry[12]), .sum(sum[14]), .cout(halfcarry[13]));
   fullAdder__0_258 genblk2_14_f3 (.x(halfsum[15]), .y(halfcout[14]), .cin(
      halfcarry[13]), .sum(sum[15]), .cout(halfcarry[14]));
   fullAdder__0_255 genblk2_15_f3 (.x(halfsum[16]), .y(halfcout[15]), .cin(
      halfcarry[14]), .sum(sum[16]), .cout(halfcarry[15]));
   fullAdder__0_252 genblk2_16_f3 (.x(halfsum[17]), .y(halfcout[16]), .cin(
      halfcarry[15]), .sum(sum[17]), .cout(halfcarry[16]));
   fullAdder__0_249 genblk2_17_f3 (.x(halfsum[18]), .y(halfcout[17]), .cin(
      halfcarry[16]), .sum(sum[18]), .cout(halfcarry[17]));
   fullAdder__0_246 genblk2_18_f3 (.x(halfsum[19]), .y(halfcout[18]), .cin(
      halfcarry[17]), .sum(sum[19]), .cout(halfcarry[18]));
   fullAdder__0_243 genblk2_19_f3 (.x(halfsum[20]), .y(halfcout[19]), .cin(
      halfcarry[18]), .sum(sum[20]), .cout(halfcarry[19]));
   fullAdder__0_240 genblk2_20_f3 (.x(halfsum[21]), .y(halfcout[20]), .cin(
      halfcarry[19]), .sum(sum[21]), .cout(halfcarry[20]));
   fullAdder__0_237 genblk2_21_f3 (.x(halfsum[22]), .y(halfcout[21]), .cin(
      halfcarry[20]), .sum(sum[22]), .cout(halfcarry[21]));
   fullAdder__0_234 genblk2_22_f3 (.x(halfsum[23]), .y(halfcout[22]), .cin(
      halfcarry[21]), .sum(sum[23]), .cout(halfcarry[22]));
   fullAdder__0_231 genblk2_23_f3 (.x(halfsum[24]), .y(halfcout[23]), .cin(
      halfcarry[22]), .sum(sum[24]), .cout(halfcarry[23]));
   fullAdder__0_228 genblk2_24_f3 (.x(halfsum[25]), .y(halfcout[24]), .cin(
      halfcarry[23]), .sum(sum[25]), .cout(halfcarry[24]));
   fullAdder__0_225 genblk2_25_f3 (.x(halfsum[26]), .y(halfcout[25]), .cin(
      halfcarry[24]), .sum(sum[26]), .cout(halfcarry[25]));
   fullAdder__0_222 genblk2_26_f3 (.x(halfsum[27]), .y(halfcout[26]), .cin(
      halfcarry[25]), .sum(sum[27]), .cout(halfcarry[26]));
   fullAdder__0_219 genblk2_27_f3 (.x(halfsum[28]), .y(halfcout[27]), .cin(
      halfcarry[26]), .sum(sum[28]), .cout(halfcarry[27]));
   fullAdder__0_216 genblk2_28_f3 (.x(halfsum[29]), .y(halfcout[28]), .cin(
      halfcarry[27]), .sum(sum[29]), .cout(halfcarry[28]));
   fullAdder__0_213 genblk2_29_f3 (.x(halfsum[30]), .y(halfcout[29]), .cin(
      halfcarry[28]), .sum(sum[30]), .cout(halfcarry[29]));
   fullAdder__0_210 genblk2_30_f3 (.x(halfsum[31]), .y(halfcout[30]), .cin(
      halfcarry[29]), .sum(sum[31]), .cout());
endmodule

module fullAdder__0_21(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_27(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_30(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_33(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_36(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_39(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_42(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_45(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_48(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_51(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_54(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_57(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_60(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_63(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_66(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_69(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_72(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_75(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_78(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_81(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_84(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_87(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_90(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_93(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_96(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_99(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_102(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_105(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_108(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_111(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_114(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_117(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_120(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(y), .B(x), .Z(sum));
endmodule

module fullAdder__0_123(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_126(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_129(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_132(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_135(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_138(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_141(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_144(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_147(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_150(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_153(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_156(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_159(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_162(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_165(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_168(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_171(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_174(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_177(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_180(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_183(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_186(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_189(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_192(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_195(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_198(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_201(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_204(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_207(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(x), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(y), .ZN(sum));
endmodule

module carrySaveAdder(a, b, c, sum, cout);
   input [31:0]a;
   input [31:0]b;
   input [31:0]c;
   output [31:0]sum;
   output cout;

   wire [31:0]halfcarry;
   wire [31:0]halfcout;
   wire [31:0]halfsum;

   fullAdder__0_21 fulladder_f2 (.x(halfsum[1]), .y(halfcout[0]), .cin(), 
      .sum(sum[1]), .cout(halfcarry[0]));
   fullAdder__0_27 genblk1_0_fulladder_f1 (.x(a[0]), .y(b[0]), .cin(), .sum(
      sum[0]), .cout(halfcout[0]));
   fullAdder__0_30 genblk1_1_fulladder_f1 (.x(a[1]), .y(b[1]), .cin(), .sum(
      halfsum[1]), .cout(halfcout[1]));
   fullAdder__0_33 genblk1_2_fulladder_f1 (.x(a[2]), .y(b[2]), .cin(), .sum(
      halfsum[2]), .cout(halfcout[2]));
   fullAdder__0_36 genblk1_3_fulladder_f1 (.x(a[3]), .y(b[3]), .cin(), .sum(
      halfsum[3]), .cout(halfcout[3]));
   fullAdder__0_39 genblk1_4_fulladder_f1 (.x(a[4]), .y(b[4]), .cin(), .sum(
      halfsum[4]), .cout(halfcout[4]));
   fullAdder__0_42 genblk1_5_fulladder_f1 (.x(a[5]), .y(b[5]), .cin(), .sum(
      halfsum[5]), .cout(halfcout[5]));
   fullAdder__0_45 genblk1_6_fulladder_f1 (.x(a[6]), .y(b[6]), .cin(), .sum(
      halfsum[6]), .cout(halfcout[6]));
   fullAdder__0_48 genblk1_7_fulladder_f1 (.x(a[7]), .y(b[7]), .cin(), .sum(
      halfsum[7]), .cout(halfcout[7]));
   fullAdder__0_51 genblk1_8_fulladder_f1 (.x(a[8]), .y(b[8]), .cin(), .sum(
      halfsum[8]), .cout(halfcout[8]));
   fullAdder__0_54 genblk1_9_fulladder_f1 (.x(a[9]), .y(b[9]), .cin(), .sum(
      halfsum[9]), .cout(halfcout[9]));
   fullAdder__0_57 genblk1_10_fulladder_f1 (.x(a[10]), .y(b[10]), .cin(), 
      .sum(halfsum[10]), .cout(halfcout[10]));
   fullAdder__0_60 genblk1_11_fulladder_f1 (.x(a[11]), .y(b[11]), .cin(), 
      .sum(halfsum[11]), .cout(halfcout[11]));
   fullAdder__0_63 genblk1_12_fulladder_f1 (.x(a[12]), .y(b[12]), .cin(), 
      .sum(halfsum[12]), .cout(halfcout[12]));
   fullAdder__0_66 genblk1_13_fulladder_f1 (.x(a[13]), .y(b[13]), .cin(), 
      .sum(halfsum[13]), .cout(halfcout[13]));
   fullAdder__0_69 genblk1_14_fulladder_f1 (.x(a[14]), .y(b[14]), .cin(), 
      .sum(halfsum[14]), .cout(halfcout[14]));
   fullAdder__0_72 genblk1_15_fulladder_f1 (.x(a[15]), .y(b[15]), .cin(), 
      .sum(halfsum[15]), .cout(halfcout[15]));
   fullAdder__0_75 genblk1_16_fulladder_f1 (.x(a[16]), .y(b[16]), .cin(), 
      .sum(halfsum[16]), .cout(halfcout[16]));
   fullAdder__0_78 genblk1_17_fulladder_f1 (.x(a[17]), .y(b[17]), .cin(), 
      .sum(halfsum[17]), .cout(halfcout[17]));
   fullAdder__0_81 genblk1_18_fulladder_f1 (.x(a[18]), .y(b[18]), .cin(), 
      .sum(halfsum[18]), .cout(halfcout[18]));
   fullAdder__0_84 genblk1_19_fulladder_f1 (.x(a[19]), .y(b[19]), .cin(), 
      .sum(halfsum[19]), .cout(halfcout[19]));
   fullAdder__0_87 genblk1_20_fulladder_f1 (.x(a[20]), .y(b[20]), .cin(), 
      .sum(halfsum[20]), .cout(halfcout[20]));
   fullAdder__0_90 genblk1_21_fulladder_f1 (.x(a[21]), .y(b[21]), .cin(), 
      .sum(halfsum[21]), .cout(halfcout[21]));
   fullAdder__0_93 genblk1_22_fulladder_f1 (.x(a[22]), .y(b[22]), .cin(), 
      .sum(halfsum[22]), .cout(halfcout[22]));
   fullAdder__0_96 genblk1_23_fulladder_f1 (.x(a[23]), .y(b[23]), .cin(), 
      .sum(halfsum[23]), .cout(halfcout[23]));
   fullAdder__0_99 genblk1_24_fulladder_f1 (.x(a[24]), .y(b[24]), .cin(), 
      .sum(halfsum[24]), .cout(halfcout[24]));
   fullAdder__0_102 genblk1_25_fulladder_f1 (.x(a[25]), .y(b[25]), .cin(), 
      .sum(halfsum[25]), .cout(halfcout[25]));
   fullAdder__0_105 genblk1_26_fulladder_f1 (.x(a[26]), .y(b[26]), .cin(), 
      .sum(halfsum[26]), .cout(halfcout[26]));
   fullAdder__0_108 genblk1_27_fulladder_f1 (.x(a[27]), .y(b[27]), .cin(), 
      .sum(halfsum[27]), .cout(halfcout[27]));
   fullAdder__0_111 genblk1_28_fulladder_f1 (.x(a[28]), .y(b[28]), .cin(), 
      .sum(halfsum[28]), .cout(halfcout[28]));
   fullAdder__0_114 genblk1_29_fulladder_f1 (.x(a[29]), .y(b[29]), .cin(), 
      .sum(halfsum[29]), .cout(halfcout[29]));
   fullAdder__0_117 genblk1_30_fulladder_f1 (.x(a[30]), .y(b[30]), .cin(), 
      .sum(halfsum[30]), .cout(halfcout[30]));
   fullAdder__0_120 genblk1_31_fulladder_f1 (.x(a[31]), .y(b[31]), .cin(), 
      .sum(halfsum[31]), .cout());
   fullAdder__0_123 genblk2_1_f3 (.x(halfsum[2]), .y(halfcout[1]), .cin(
      halfcarry[0]), .sum(sum[2]), .cout(halfcarry[1]));
   fullAdder__0_126 genblk2_2_f3 (.x(halfsum[3]), .y(halfcout[2]), .cin(
      halfcarry[1]), .sum(sum[3]), .cout(halfcarry[2]));
   fullAdder__0_129 genblk2_3_f3 (.x(halfsum[4]), .y(halfcout[3]), .cin(
      halfcarry[2]), .sum(sum[4]), .cout(halfcarry[3]));
   fullAdder__0_132 genblk2_4_f3 (.x(halfsum[5]), .y(halfcout[4]), .cin(
      halfcarry[3]), .sum(sum[5]), .cout(halfcarry[4]));
   fullAdder__0_135 genblk2_5_f3 (.x(halfsum[6]), .y(halfcout[5]), .cin(
      halfcarry[4]), .sum(sum[6]), .cout(halfcarry[5]));
   fullAdder__0_138 genblk2_6_f3 (.x(halfsum[7]), .y(halfcout[6]), .cin(
      halfcarry[5]), .sum(sum[7]), .cout(halfcarry[6]));
   fullAdder__0_141 genblk2_7_f3 (.x(halfsum[8]), .y(halfcout[7]), .cin(
      halfcarry[6]), .sum(sum[8]), .cout(halfcarry[7]));
   fullAdder__0_144 genblk2_8_f3 (.x(halfsum[9]), .y(halfcout[8]), .cin(
      halfcarry[7]), .sum(sum[9]), .cout(halfcarry[8]));
   fullAdder__0_147 genblk2_9_f3 (.x(halfsum[10]), .y(halfcout[9]), .cin(
      halfcarry[8]), .sum(sum[10]), .cout(halfcarry[9]));
   fullAdder__0_150 genblk2_10_f3 (.x(halfsum[11]), .y(halfcout[10]), .cin(
      halfcarry[9]), .sum(sum[11]), .cout(halfcarry[10]));
   fullAdder__0_153 genblk2_11_f3 (.x(halfsum[12]), .y(halfcout[11]), .cin(
      halfcarry[10]), .sum(sum[12]), .cout(halfcarry[11]));
   fullAdder__0_156 genblk2_12_f3 (.x(halfsum[13]), .y(halfcout[12]), .cin(
      halfcarry[11]), .sum(sum[13]), .cout(halfcarry[12]));
   fullAdder__0_159 genblk2_13_f3 (.x(halfsum[14]), .y(halfcout[13]), .cin(
      halfcarry[12]), .sum(sum[14]), .cout(halfcarry[13]));
   fullAdder__0_162 genblk2_14_f3 (.x(halfsum[15]), .y(halfcout[14]), .cin(
      halfcarry[13]), .sum(sum[15]), .cout(halfcarry[14]));
   fullAdder__0_165 genblk2_15_f3 (.x(halfsum[16]), .y(halfcout[15]), .cin(
      halfcarry[14]), .sum(sum[16]), .cout(halfcarry[15]));
   fullAdder__0_168 genblk2_16_f3 (.x(halfsum[17]), .y(halfcout[16]), .cin(
      halfcarry[15]), .sum(sum[17]), .cout(halfcarry[16]));
   fullAdder__0_171 genblk2_17_f3 (.x(halfsum[18]), .y(halfcout[17]), .cin(
      halfcarry[16]), .sum(sum[18]), .cout(halfcarry[17]));
   fullAdder__0_174 genblk2_18_f3 (.x(halfsum[19]), .y(halfcout[18]), .cin(
      halfcarry[17]), .sum(sum[19]), .cout(halfcarry[18]));
   fullAdder__0_177 genblk2_19_f3 (.x(halfsum[20]), .y(halfcout[19]), .cin(
      halfcarry[18]), .sum(sum[20]), .cout(halfcarry[19]));
   fullAdder__0_180 genblk2_20_f3 (.x(halfsum[21]), .y(halfcout[20]), .cin(
      halfcarry[19]), .sum(sum[21]), .cout(halfcarry[20]));
   fullAdder__0_183 genblk2_21_f3 (.x(halfsum[22]), .y(halfcout[21]), .cin(
      halfcarry[20]), .sum(sum[22]), .cout(halfcarry[21]));
   fullAdder__0_186 genblk2_22_f3 (.x(halfsum[23]), .y(halfcout[22]), .cin(
      halfcarry[21]), .sum(sum[23]), .cout(halfcarry[22]));
   fullAdder__0_189 genblk2_23_f3 (.x(halfsum[24]), .y(halfcout[23]), .cin(
      halfcarry[22]), .sum(sum[24]), .cout(halfcarry[23]));
   fullAdder__0_192 genblk2_24_f3 (.x(halfsum[25]), .y(halfcout[24]), .cin(
      halfcarry[23]), .sum(sum[25]), .cout(halfcarry[24]));
   fullAdder__0_195 genblk2_25_f3 (.x(halfsum[26]), .y(halfcout[25]), .cin(
      halfcarry[24]), .sum(sum[26]), .cout(halfcarry[25]));
   fullAdder__0_198 genblk2_26_f3 (.x(halfsum[27]), .y(halfcout[26]), .cin(
      halfcarry[25]), .sum(sum[27]), .cout(halfcarry[26]));
   fullAdder__0_201 genblk2_27_f3 (.x(halfsum[28]), .y(halfcout[27]), .cin(
      halfcarry[26]), .sum(sum[28]), .cout(halfcarry[27]));
   fullAdder__0_204 genblk2_28_f3 (.x(halfsum[29]), .y(halfcout[28]), .cin(
      halfcarry[27]), .sum(sum[29]), .cout(halfcarry[28]));
   fullAdder__0_207 genblk2_29_f3 (.x(halfsum[30]), .y(halfcout[29]), .cin(
      halfcarry[28]), .sum(sum[30]), .cout(halfcarry[29]));
   fullAdder genblk2_30_f3 (.x(halfsum[31]), .y(halfcout[30]), .cin(
      halfcarry[29]), .sum(sum[31]), .cout());
endmodule

module regFile(read_data, read_data2, write_en, write_data, write_data2, clk);
   output [31:0]read_data;
   output [31:0]read_data2;
   input write_en;
   input [31:0]write_data;
   input [31:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[31]  (.D(write_data2[31]), .CK(n_0), .Q(read_data2[31]), 
      .QN());
   DFF_X1 \my_reg2_reg[30]  (.D(write_data2[30]), .CK(n_0), .Q(read_data2[30]), 
      .QN());
   DFF_X1 \my_reg2_reg[29]  (.D(write_data2[29]), .CK(n_0), .Q(read_data2[29]), 
      .QN());
   DFF_X1 \my_reg2_reg[28]  (.D(write_data2[28]), .CK(n_0), .Q(read_data2[28]), 
      .QN());
   DFF_X1 \my_reg2_reg[27]  (.D(write_data2[27]), .CK(n_0), .Q(read_data2[27]), 
      .QN());
   DFF_X1 \my_reg2_reg[26]  (.D(write_data2[26]), .CK(n_0), .Q(read_data2[26]), 
      .QN());
   DFF_X1 \my_reg2_reg[25]  (.D(write_data2[25]), .CK(n_0), .Q(read_data2[25]), 
      .QN());
   DFF_X1 \my_reg2_reg[24]  (.D(write_data2[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data2[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
   DFF_X1 \my_reg2_reg[22]  (.D(write_data2[22]), .CK(n_0), .Q(read_data2[22]), 
      .QN());
   DFF_X1 \my_reg2_reg[21]  (.D(write_data2[21]), .CK(n_0), .Q(read_data2[21]), 
      .QN());
   DFF_X1 \my_reg2_reg[20]  (.D(write_data2[20]), .CK(n_0), .Q(read_data2[20]), 
      .QN());
   DFF_X1 \my_reg2_reg[19]  (.D(write_data2[19]), .CK(n_0), .Q(read_data2[19]), 
      .QN());
   DFF_X1 \my_reg2_reg[18]  (.D(write_data2[18]), .CK(n_0), .Q(read_data2[18]), 
      .QN());
   DFF_X1 \my_reg2_reg[17]  (.D(write_data2[17]), .CK(n_0), .Q(read_data2[17]), 
      .QN());
   DFF_X1 \my_reg2_reg[16]  (.D(write_data2[16]), .CK(n_0), .Q(read_data2[16]), 
      .QN());
   DFF_X1 \my_reg2_reg[15]  (.D(write_data2[15]), .CK(n_0), .Q(read_data2[15]), 
      .QN());
   DFF_X1 \my_reg2_reg[14]  (.D(write_data2[14]), .CK(n_0), .Q(read_data2[14]), 
      .QN());
   DFF_X1 \my_reg2_reg[13]  (.D(write_data2[13]), .CK(n_0), .Q(read_data2[13]), 
      .QN());
   DFF_X1 \my_reg2_reg[12]  (.D(write_data2[12]), .CK(n_0), .Q(read_data2[12]), 
      .QN());
   DFF_X1 \my_reg2_reg[11]  (.D(write_data2[11]), .CK(n_0), .Q(read_data2[11]), 
      .QN());
   DFF_X1 \my_reg2_reg[10]  (.D(write_data2[10]), .CK(n_0), .Q(read_data2[10]), 
      .QN());
   DFF_X1 \my_reg2_reg[9]  (.D(write_data2[9]), .CK(n_0), .Q(read_data2[9]), 
      .QN());
   DFF_X1 \my_reg2_reg[8]  (.D(write_data2[8]), .CK(n_0), .Q(read_data2[8]), 
      .QN());
   DFF_X1 \my_reg2_reg[7]  (.D(write_data2[7]), .CK(n_0), .Q(read_data2[7]), 
      .QN());
   DFF_X1 \my_reg2_reg[6]  (.D(write_data2[6]), .CK(n_0), .Q(read_data2[6]), 
      .QN());
   DFF_X1 \my_reg2_reg[5]  (.D(write_data2[5]), .CK(n_0), .Q(read_data2[5]), 
      .QN());
   DFF_X1 \my_reg2_reg[4]  (.D(write_data2[4]), .CK(n_0), .Q(read_data2[4]), 
      .QN());
   DFF_X1 \my_reg2_reg[3]  (.D(write_data2[3]), .CK(n_0), .Q(read_data2[3]), 
      .QN());
   DFF_X1 \my_reg2_reg[2]  (.D(write_data2[2]), .CK(n_0), .Q(read_data2[2]), 
      .QN());
   DFF_X1 \my_reg2_reg[1]  (.D(write_data2[1]), .CK(n_0), .Q(read_data2[1]), 
      .QN());
   DFF_X1 \my_reg2_reg[0]  (.D(write_data2[0]), .CK(n_0), .Q(read_data2[0]), 
      .QN());
   DFF_X1 \my_reg_reg[31]  (.D(write_data[31]), .CK(n_0), .Q(read_data[31]), 
      .QN());
   DFF_X1 \my_reg_reg[30]  (.D(write_data[30]), .CK(n_0), .Q(read_data[30]), 
      .QN());
   DFF_X1 \my_reg_reg[29]  (.D(write_data[29]), .CK(n_0), .Q(read_data[29]), 
      .QN());
   DFF_X1 \my_reg_reg[28]  (.D(write_data[28]), .CK(n_0), .Q(read_data[28]), 
      .QN());
   DFF_X1 \my_reg_reg[27]  (.D(write_data[27]), .CK(n_0), .Q(read_data[27]), 
      .QN());
   DFF_X1 \my_reg_reg[26]  (.D(write_data[26]), .CK(n_0), .Q(read_data[26]), 
      .QN());
   DFF_X1 \my_reg_reg[25]  (.D(write_data[25]), .CK(n_0), .Q(read_data[25]), 
      .QN());
   DFF_X1 \my_reg_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data[24]), 
      .QN());
   DFF_X1 \my_reg_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data[23]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
endmodule

module datapath__0_17(f8, p_0);
   input [31:0]f8;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(f8[1]), .B(f8[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(f8[2]), .B1(f8[1]), .B2(f8[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(f8[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(f8[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(f8[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(f8[6]), .B1(n_27), .B2(f8[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(f8[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(f8[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(f8[9]), .B1(n_25), .B2(f8[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(f8[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(f8[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(f8[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(f8[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(f8[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(f8[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(f8[16]), .B1(n_19), .B2(f8[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(f8[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(f8[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(f8[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(f8[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(f8[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(f8[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(f8[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(f8[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(f8[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(f8[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(f8[27]), .B1(n_9), .B2(f8[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(f8[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(f8[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(f8[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(f8[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(f8[28]), .A3(f8[29]), .A4(f8[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(f8[28]), .A3(f8[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(f8[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(f8[26]), .A3(f8[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(f8[23]), .A3(f8[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(f8[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(f8[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(f8[18]), .A3(f8[19]), .A4(f8[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(f8[18]), .A3(f8[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(f8[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(f8[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(f8[15]), .A3(f8[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(f8[12]), .A3(f8[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(f8[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(f8[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(f8[8]), .A3(f8[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(f8[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(f8[5]), .A3(f8[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(f8[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(f8[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(f8[2]), .A2(f8[1]), .A3(f8[0]), .ZN(n_29));
   INV_X1 i_61 (.A(f8[11]), .ZN(n_30));
   INV_X1 i_62 (.A(f8[14]), .ZN(n_31));
   INV_X1 i_63 (.A(f8[21]), .ZN(n_32));
   INV_X1 i_64 (.A(f8[25]), .ZN(n_33));
endmodule

module BoothAlgo(M, Q, result, clk, start);
   input [31:0]M;
   input [31:0]Q;
   output [63:0]result;
   input clk;
   input start;

   wire [31:0]read2;
   wire [31:0]read;
   wire [31:0]SubM;
   wire [31:0]AddM;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire [31:0]A;
   wire n_0_102;
   wire [31:0]l8;
   wire n_0_31;
   wire [31:0]f8;
   wire write_en;
   wire write_en2;
   wire n_0_103;
   wire [5:0]count;
   wire q0;
   wire n_0_32;
   wire n_0_34;
   wire n_0_35;
   wire n_0_1_0;
   wire n_0_36;
   wire n_0_1_1;
   wire n_0_37;
   wire n_0_1_2;
   wire n_0_38;
   wire n_0_1_3;
   wire n_0_39;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_40;
   wire n_0_41;
   wire n_0_1_8;
   wire n_0_42;
   wire n_0_1_9;
   wire n_0_43;
   wire n_0_1_10;
   wire n_0_44;
   wire n_0_1_11;
   wire n_0_45;
   wire n_0_1_12;
   wire n_0_46;
   wire n_0_1_13;
   wire n_0_47;
   wire n_0_1_14;
   wire n_0_48;
   wire n_0_1_15;
   wire n_0_49;
   wire n_0_1_16;
   wire n_0_50;
   wire n_0_1_17;
   wire n_0_51;
   wire n_0_1_18;
   wire n_0_52;
   wire n_0_1_19;
   wire n_0_53;
   wire n_0_1_20;
   wire n_0_54;
   wire n_0_1_21;
   wire n_0_55;
   wire n_0_1_22;
   wire n_0_56;
   wire n_0_1_23;
   wire n_0_57;
   wire n_0_1_24;
   wire n_0_58;
   wire n_0_1_25;
   wire n_0_59;
   wire n_0_1_26;
   wire n_0_60;
   wire n_0_1_27;
   wire n_0_61;
   wire n_0_1_28;
   wire n_0_62;
   wire n_0_1_29;
   wire n_0_63;
   wire n_0_1_30;
   wire n_0_64;
   wire n_0_1_31;
   wire n_0_65;
   wire n_0_1_32;
   wire n_0_66;
   wire n_0_1_33;
   wire n_0_67;
   wire n_0_1_34;
   wire n_0_68;
   wire n_0_1_35;
   wire n_0_69;
   wire n_0_1_36;
   wire n_0_70;
   wire n_0_1_37;
   wire n_0_71;
   wire n_0_1_38;
   wire n_0_72;
   wire n_0_1_39;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_101;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_99;
   wire n_0_100;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_33;
   wire n_0_1_49;

   regFile__0_18 inst1 (.read_data(read), .read_data2(read2), .write_en(write_en), 
      .write_data(M), .write_data2(Q), .clk(clk));
   carrySaveAdder__0_400 subtractor (.a(A), .b({n_0_30, n_0_29, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, 
      n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, f8[0]}), 
      .c(), .sum(SubM), .cout());
   carrySaveAdder adder (.a(A), .b(f8), .c(), .sum(AddM), .cout());
   regFile inst2 (.read_data({result[63], result[62], result[61], result[60], 
      result[59], result[58], result[57], result[56], result[55], result[54], 
      result[53], result[52], result[51], result[50], result[49], result[48], 
      result[47], result[46], result[45], result[44], result[43], result[42], 
      result[41], result[40], result[39], result[38], result[37], result[36], 
      result[35], result[34], result[33], result[32]}), .read_data2({result[31], 
      result[30], result[29], result[28], result[27], result[26], result[25], 
      result[24], result[23], result[22], result[21], result[20], result[19], 
      result[18], result[17], result[16], result[15], result[14], result[13], 
      result[12], result[11], result[10], result[9], result[8], result[7], 
      result[6], result[5], result[4], result[3], result[2], result[1], 
      result[0]}), .write_en(write_en2), .write_data(A), .write_data2(l8), 
      .clk(clk));
   datapath__0_17 i_0_0 (.f8(f8), .p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_0}));
   DFF_X1 \A_reg[30]  (.D(n_0_71), .CK(n_0_32), .Q(A[30]), .QN());
   DFF_X1 \A_reg[29]  (.D(n_0_70), .CK(n_0_32), .Q(A[29]), .QN());
   DFF_X1 \A_reg[28]  (.D(n_0_69), .CK(n_0_32), .Q(A[28]), .QN());
   DFF_X1 \A_reg[27]  (.D(n_0_68), .CK(n_0_32), .Q(A[27]), .QN());
   DFF_X1 \A_reg[26]  (.D(n_0_67), .CK(n_0_32), .Q(A[26]), .QN());
   DFF_X1 \A_reg[25]  (.D(n_0_66), .CK(n_0_32), .Q(A[25]), .QN());
   DFF_X1 \A_reg[24]  (.D(n_0_65), .CK(n_0_32), .Q(A[24]), .QN());
   DFF_X1 \A_reg[23]  (.D(n_0_64), .CK(n_0_32), .Q(A[23]), .QN());
   DFF_X1 \A_reg[22]  (.D(n_0_63), .CK(n_0_32), .Q(A[22]), .QN());
   DFF_X1 \A_reg[21]  (.D(n_0_62), .CK(n_0_32), .Q(A[21]), .QN());
   DFF_X1 \A_reg[20]  (.D(n_0_61), .CK(n_0_32), .Q(A[20]), .QN());
   DFF_X1 \A_reg[19]  (.D(n_0_60), .CK(n_0_32), .Q(A[19]), .QN());
   DFF_X1 \A_reg[18]  (.D(n_0_59), .CK(n_0_32), .Q(A[18]), .QN());
   DFF_X1 \A_reg[17]  (.D(n_0_58), .CK(n_0_32), .Q(A[17]), .QN());
   DFF_X1 \A_reg[16]  (.D(n_0_57), .CK(n_0_32), .Q(A[16]), .QN());
   DFF_X1 \A_reg[15]  (.D(n_0_56), .CK(n_0_32), .Q(A[15]), .QN());
   DFF_X1 \A_reg[14]  (.D(n_0_55), .CK(n_0_32), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(n_0_54), .CK(n_0_32), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(n_0_53), .CK(n_0_32), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(n_0_52), .CK(n_0_32), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(n_0_51), .CK(n_0_32), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(n_0_50), .CK(n_0_32), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(n_0_49), .CK(n_0_32), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(n_0_48), .CK(n_0_32), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(n_0_47), .CK(n_0_32), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(n_0_46), .CK(n_0_32), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(n_0_45), .CK(n_0_32), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(n_0_44), .CK(n_0_32), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(n_0_43), .CK(n_0_32), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(n_0_42), .CK(n_0_32), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(n_0_41), .CK(n_0_32), .Q(A[0]), .QN());
   DFF_X1 \A_reg[31]  (.D(n_0_102), .CK(clk), .Q(A[31]), .QN());
   MUX2_X1 \A_reg[31]_enable_mux_0  (.A(A[31]), .B(n_0_72), .S(n_0_101), 
      .Z(n_0_102));
   DFF_X1 \l8_reg[31]  (.D(n_0_98), .CK(n_0_32), .Q(l8[31]), .QN());
   DFF_X1 \l8_reg[30]  (.D(n_0_97), .CK(n_0_32), .Q(l8[30]), .QN());
   DFF_X1 \l8_reg[29]  (.D(n_0_96), .CK(n_0_32), .Q(l8[29]), .QN());
   DFF_X1 \l8_reg[28]  (.D(n_0_95), .CK(n_0_32), .Q(l8[28]), .QN());
   DFF_X1 \l8_reg[27]  (.D(n_0_94), .CK(n_0_32), .Q(l8[27]), .QN());
   DFF_X1 \l8_reg[26]  (.D(n_0_93), .CK(n_0_32), .Q(l8[26]), .QN());
   DFF_X1 \l8_reg[25]  (.D(n_0_92), .CK(n_0_32), .Q(l8[25]), .QN());
   DFF_X1 \l8_reg[24]  (.D(n_0_91), .CK(n_0_32), .Q(l8[24]), .QN());
   DFF_X1 \l8_reg[23]  (.D(n_0_90), .CK(n_0_32), .Q(l8[23]), .QN());
   DFF_X1 \l8_reg[22]  (.D(n_0_89), .CK(n_0_32), .Q(l8[22]), .QN());
   DFF_X1 \l8_reg[21]  (.D(n_0_88), .CK(n_0_32), .Q(l8[21]), .QN());
   DFF_X1 \l8_reg[20]  (.D(n_0_87), .CK(n_0_32), .Q(l8[20]), .QN());
   DFF_X1 \l8_reg[19]  (.D(n_0_86), .CK(n_0_32), .Q(l8[19]), .QN());
   DFF_X1 \l8_reg[18]  (.D(n_0_85), .CK(n_0_32), .Q(l8[18]), .QN());
   DFF_X1 \l8_reg[17]  (.D(n_0_84), .CK(n_0_32), .Q(l8[17]), .QN());
   DFF_X1 \l8_reg[16]  (.D(n_0_83), .CK(n_0_32), .Q(l8[16]), .QN());
   DFF_X1 \l8_reg[15]  (.D(n_0_82), .CK(n_0_32), .Q(l8[15]), .QN());
   DFF_X1 \l8_reg[14]  (.D(n_0_81), .CK(n_0_32), .Q(l8[14]), .QN());
   DFF_X1 \l8_reg[13]  (.D(n_0_80), .CK(n_0_32), .Q(l8[13]), .QN());
   DFF_X1 \l8_reg[12]  (.D(n_0_79), .CK(n_0_32), .Q(l8[12]), .QN());
   DFF_X1 \l8_reg[11]  (.D(n_0_78), .CK(n_0_32), .Q(l8[11]), .QN());
   DFF_X1 \l8_reg[10]  (.D(n_0_77), .CK(n_0_32), .Q(l8[10]), .QN());
   DFF_X1 \l8_reg[9]  (.D(n_0_76), .CK(n_0_32), .Q(l8[9]), .QN());
   DFF_X1 \l8_reg[8]  (.D(n_0_75), .CK(n_0_32), .Q(l8[8]), .QN());
   DFF_X1 \l8_reg[7]  (.D(n_0_74), .CK(n_0_32), .Q(l8[7]), .QN());
   DFF_X1 \l8_reg[6]  (.D(n_0_73), .CK(n_0_32), .Q(l8[6]), .QN());
   DFF_X1 \l8_reg[5]  (.D(n_0_109), .CK(n_0_32), .Q(l8[5]), .QN());
   DFF_X1 \l8_reg[4]  (.D(n_0_108), .CK(n_0_32), .Q(l8[4]), .QN());
   DFF_X1 \l8_reg[3]  (.D(n_0_107), .CK(n_0_32), .Q(l8[3]), .QN());
   DFF_X1 \l8_reg[2]  (.D(n_0_106), .CK(n_0_32), .Q(l8[2]), .QN());
   DFF_X1 \l8_reg[1]  (.D(n_0_105), .CK(n_0_32), .Q(l8[1]), .QN());
   DFF_X1 \l8_reg[0]  (.D(n_0_104), .CK(n_0_32), .Q(l8[0]), .QN());
   CLKGATETST_X1 clk_gate_f8_reg (.CK(clk), .E(start), .SE(1'b0), .GCK(n_0_31));
   DFF_X1 \f8_reg[31]  (.D(read[31]), .CK(n_0_31), .Q(f8[31]), .QN());
   DFF_X1 \f8_reg[30]  (.D(read[30]), .CK(n_0_31), .Q(f8[30]), .QN());
   DFF_X1 \f8_reg[29]  (.D(read[29]), .CK(n_0_31), .Q(f8[29]), .QN());
   DFF_X1 \f8_reg[28]  (.D(read[28]), .CK(n_0_31), .Q(f8[28]), .QN());
   DFF_X1 \f8_reg[27]  (.D(read[27]), .CK(n_0_31), .Q(f8[27]), .QN());
   DFF_X1 \f8_reg[26]  (.D(read[26]), .CK(n_0_31), .Q(f8[26]), .QN());
   DFF_X1 \f8_reg[25]  (.D(read[25]), .CK(n_0_31), .Q(f8[25]), .QN());
   DFF_X1 \f8_reg[24]  (.D(read[24]), .CK(n_0_31), .Q(f8[24]), .QN());
   DFF_X1 \f8_reg[23]  (.D(read[23]), .CK(n_0_31), .Q(f8[23]), .QN());
   DFF_X1 \f8_reg[22]  (.D(read[22]), .CK(n_0_31), .Q(f8[22]), .QN());
   DFF_X1 \f8_reg[21]  (.D(read[21]), .CK(n_0_31), .Q(f8[21]), .QN());
   DFF_X1 \f8_reg[20]  (.D(read[20]), .CK(n_0_31), .Q(f8[20]), .QN());
   DFF_X1 \f8_reg[19]  (.D(read[19]), .CK(n_0_31), .Q(f8[19]), .QN());
   DFF_X1 \f8_reg[18]  (.D(read[18]), .CK(n_0_31), .Q(f8[18]), .QN());
   DFF_X1 \f8_reg[17]  (.D(read[17]), .CK(n_0_31), .Q(f8[17]), .QN());
   DFF_X1 \f8_reg[16]  (.D(read[16]), .CK(n_0_31), .Q(f8[16]), .QN());
   DFF_X1 \f8_reg[15]  (.D(read[15]), .CK(n_0_31), .Q(f8[15]), .QN());
   DFF_X1 \f8_reg[14]  (.D(read[14]), .CK(n_0_31), .Q(f8[14]), .QN());
   DFF_X1 \f8_reg[13]  (.D(read[13]), .CK(n_0_31), .Q(f8[13]), .QN());
   DFF_X1 \f8_reg[12]  (.D(read[12]), .CK(n_0_31), .Q(f8[12]), .QN());
   DFF_X1 \f8_reg[11]  (.D(read[11]), .CK(n_0_31), .Q(f8[11]), .QN());
   DFF_X1 \f8_reg[10]  (.D(read[10]), .CK(n_0_31), .Q(f8[10]), .QN());
   DFF_X1 \f8_reg[9]  (.D(read[9]), .CK(n_0_31), .Q(f8[9]), .QN());
   DFF_X1 \f8_reg[8]  (.D(read[8]), .CK(n_0_31), .Q(f8[8]), .QN());
   DFF_X1 \f8_reg[7]  (.D(read[7]), .CK(n_0_31), .Q(f8[7]), .QN());
   DFF_X1 \f8_reg[6]  (.D(read[6]), .CK(n_0_31), .Q(f8[6]), .QN());
   DFF_X1 \f8_reg[5]  (.D(read[5]), .CK(n_0_31), .Q(f8[5]), .QN());
   DFF_X1 \f8_reg[4]  (.D(read[4]), .CK(n_0_31), .Q(f8[4]), .QN());
   DFF_X1 \f8_reg[3]  (.D(read[3]), .CK(n_0_31), .Q(f8[3]), .QN());
   DFF_X1 \f8_reg[2]  (.D(read[2]), .CK(n_0_31), .Q(f8[2]), .QN());
   DFF_X1 \f8_reg[1]  (.D(read[1]), .CK(n_0_31), .Q(f8[1]), .QN());
   DFF_X1 \f8_reg[0]  (.D(read[0]), .CK(n_0_31), .Q(f8[0]), .QN());
   DFF_X1 write_en_reg (.D(start), .CK(clk), .Q(write_en), .QN());
   DFF_X1 write_en2_reg (.D(n_0_103), .CK(clk), .Q(write_en2), .QN());
   MUX2_X1 write_en2_reg_enable_mux_0 (.A(write_en2), .B(n_0_33), .S(n_0_40), 
      .Z(n_0_103));
   DFF_X1 \count_reg[5]  (.D(n_0_39), .CK(n_0_32), .Q(count[5]), .QN());
   DFF_X1 \count_reg[4]  (.D(n_0_38), .CK(n_0_32), .Q(count[4]), .QN());
   DFF_X1 \count_reg[3]  (.D(n_0_37), .CK(n_0_32), .Q(count[3]), .QN());
   DFF_X1 \count_reg[2]  (.D(n_0_36), .CK(n_0_32), .Q(count[2]), .QN());
   DFF_X1 \count_reg[1]  (.D(n_0_35), .CK(n_0_32), .Q(count[1]), .QN());
   DFF_X1 \count_reg[0]  (.D(n_0_34), .CK(n_0_32), .Q(count[0]), .QN());
   DFF_X1 q0_reg (.D(n_0_99), .CK(n_0_32), .Q(q0), .QN());
   CLKGATETST_X1 clk_gate_A_reg__0 (.CK(clk), .E(n_0_100), .SE(1'b0), .GCK(
      n_0_32));
   NOR2_X1 i_0_1_0 (.A1(start), .A2(count[0]), .ZN(n_0_34));
   AOI21_X1 i_0_1_1 (.A(n_0_1_0), .B1(count[0]), .B2(count[1]), .ZN(n_0_35));
   OAI21_X1 i_0_1_2 (.A(n_0_33), .B1(count[1]), .B2(count[0]), .ZN(n_0_1_0));
   NOR3_X1 i_0_1_3 (.A1(start), .A2(n_0_1_7), .A3(n_0_1_1), .ZN(n_0_36));
   AOI21_X1 i_0_1_4 (.A(count[2]), .B1(count[1]), .B2(count[0]), .ZN(n_0_1_1));
   NOR2_X1 i_0_1_5 (.A1(n_0_1_6), .A2(n_0_1_2), .ZN(n_0_37));
   OAI21_X1 i_0_1_6 (.A(n_0_33), .B1(count[3]), .B2(n_0_1_7), .ZN(n_0_1_2));
   NOR2_X1 i_0_1_7 (.A1(n_0_1_5), .A2(n_0_1_3), .ZN(n_0_38));
   OAI21_X1 i_0_1_8 (.A(n_0_33), .B1(count[4]), .B2(n_0_1_6), .ZN(n_0_1_3));
   NOR2_X1 i_0_1_9 (.A1(start), .A2(n_0_1_4), .ZN(n_0_39));
   XNOR2_X1 i_0_1_10 (.A(count[5]), .B(n_0_1_5), .ZN(n_0_1_4));
   AND2_X1 i_0_1_11 (.A1(count[4]), .A2(n_0_1_6), .ZN(n_0_1_5));
   AND2_X1 i_0_1_12 (.A1(count[3]), .A2(n_0_1_7), .ZN(n_0_1_6));
   AND3_X1 i_0_1_13 (.A1(count[2]), .A2(count[1]), .A3(count[0]), .ZN(n_0_1_7));
   OR2_X1 i_0_1_14 (.A1(start), .A2(n_0_1_46), .ZN(n_0_40));
   INV_X1 i_0_1_15 (.A(n_0_1_8), .ZN(n_0_41));
   AOI222_X1 i_0_1_16 (.A1(n_0_1_44), .A2(A[1]), .B1(SubM[1]), .B2(n_0_1_42), 
      .C1(AddM[1]), .C2(n_0_1_43), .ZN(n_0_1_8));
   INV_X1 i_0_1_17 (.A(n_0_1_9), .ZN(n_0_42));
   AOI222_X1 i_0_1_18 (.A1(n_0_1_44), .A2(A[2]), .B1(SubM[2]), .B2(n_0_1_42), 
      .C1(AddM[2]), .C2(n_0_1_43), .ZN(n_0_1_9));
   INV_X1 i_0_1_19 (.A(n_0_1_10), .ZN(n_0_43));
   AOI222_X1 i_0_1_20 (.A1(n_0_1_44), .A2(A[3]), .B1(SubM[3]), .B2(n_0_1_42), 
      .C1(AddM[3]), .C2(n_0_1_43), .ZN(n_0_1_10));
   INV_X1 i_0_1_21 (.A(n_0_1_11), .ZN(n_0_44));
   AOI222_X1 i_0_1_22 (.A1(n_0_1_44), .A2(A[4]), .B1(SubM[4]), .B2(n_0_1_42), 
      .C1(AddM[4]), .C2(n_0_1_43), .ZN(n_0_1_11));
   INV_X1 i_0_1_23 (.A(n_0_1_12), .ZN(n_0_45));
   AOI222_X1 i_0_1_24 (.A1(n_0_1_44), .A2(A[5]), .B1(SubM[5]), .B2(n_0_1_42), 
      .C1(AddM[5]), .C2(n_0_1_43), .ZN(n_0_1_12));
   INV_X1 i_0_1_25 (.A(n_0_1_13), .ZN(n_0_46));
   AOI222_X1 i_0_1_26 (.A1(n_0_1_44), .A2(A[6]), .B1(SubM[6]), .B2(n_0_1_42), 
      .C1(AddM[6]), .C2(n_0_1_43), .ZN(n_0_1_13));
   INV_X1 i_0_1_27 (.A(n_0_1_14), .ZN(n_0_47));
   AOI222_X1 i_0_1_28 (.A1(n_0_1_44), .A2(A[7]), .B1(SubM[7]), .B2(n_0_1_42), 
      .C1(AddM[7]), .C2(n_0_1_43), .ZN(n_0_1_14));
   INV_X1 i_0_1_29 (.A(n_0_1_15), .ZN(n_0_48));
   AOI222_X1 i_0_1_30 (.A1(n_0_1_44), .A2(A[8]), .B1(SubM[8]), .B2(n_0_1_42), 
      .C1(AddM[8]), .C2(n_0_1_43), .ZN(n_0_1_15));
   INV_X1 i_0_1_31 (.A(n_0_1_16), .ZN(n_0_49));
   AOI222_X1 i_0_1_32 (.A1(n_0_1_44), .A2(A[9]), .B1(SubM[9]), .B2(n_0_1_42), 
      .C1(AddM[9]), .C2(n_0_1_43), .ZN(n_0_1_16));
   INV_X1 i_0_1_33 (.A(n_0_1_17), .ZN(n_0_50));
   AOI222_X1 i_0_1_34 (.A1(n_0_1_44), .A2(A[10]), .B1(SubM[10]), .B2(n_0_1_42), 
      .C1(AddM[10]), .C2(n_0_1_43), .ZN(n_0_1_17));
   INV_X1 i_0_1_35 (.A(n_0_1_18), .ZN(n_0_51));
   AOI222_X1 i_0_1_36 (.A1(n_0_1_44), .A2(A[11]), .B1(SubM[11]), .B2(n_0_1_42), 
      .C1(AddM[11]), .C2(n_0_1_43), .ZN(n_0_1_18));
   INV_X1 i_0_1_37 (.A(n_0_1_19), .ZN(n_0_52));
   AOI222_X1 i_0_1_38 (.A1(n_0_1_44), .A2(A[12]), .B1(SubM[12]), .B2(n_0_1_42), 
      .C1(AddM[12]), .C2(n_0_1_43), .ZN(n_0_1_19));
   INV_X1 i_0_1_39 (.A(n_0_1_20), .ZN(n_0_53));
   AOI222_X1 i_0_1_40 (.A1(n_0_1_44), .A2(A[13]), .B1(SubM[13]), .B2(n_0_1_42), 
      .C1(AddM[13]), .C2(n_0_1_43), .ZN(n_0_1_20));
   INV_X1 i_0_1_41 (.A(n_0_1_21), .ZN(n_0_54));
   AOI222_X1 i_0_1_42 (.A1(n_0_1_44), .A2(A[14]), .B1(SubM[14]), .B2(n_0_1_42), 
      .C1(AddM[14]), .C2(n_0_1_43), .ZN(n_0_1_21));
   INV_X1 i_0_1_43 (.A(n_0_1_22), .ZN(n_0_55));
   AOI222_X1 i_0_1_44 (.A1(n_0_1_44), .A2(A[15]), .B1(SubM[15]), .B2(n_0_1_42), 
      .C1(AddM[15]), .C2(n_0_1_43), .ZN(n_0_1_22));
   INV_X1 i_0_1_45 (.A(n_0_1_23), .ZN(n_0_56));
   AOI222_X1 i_0_1_46 (.A1(n_0_1_44), .A2(A[16]), .B1(SubM[16]), .B2(n_0_1_42), 
      .C1(AddM[16]), .C2(n_0_1_43), .ZN(n_0_1_23));
   INV_X1 i_0_1_47 (.A(n_0_1_24), .ZN(n_0_57));
   AOI222_X1 i_0_1_48 (.A1(n_0_1_44), .A2(A[17]), .B1(SubM[17]), .B2(n_0_1_42), 
      .C1(AddM[17]), .C2(n_0_1_43), .ZN(n_0_1_24));
   INV_X1 i_0_1_49 (.A(n_0_1_25), .ZN(n_0_58));
   AOI222_X1 i_0_1_50 (.A1(n_0_1_44), .A2(A[18]), .B1(SubM[18]), .B2(n_0_1_42), 
      .C1(AddM[18]), .C2(n_0_1_43), .ZN(n_0_1_25));
   INV_X1 i_0_1_51 (.A(n_0_1_26), .ZN(n_0_59));
   AOI222_X1 i_0_1_52 (.A1(n_0_1_44), .A2(A[19]), .B1(SubM[19]), .B2(n_0_1_42), 
      .C1(AddM[19]), .C2(n_0_1_43), .ZN(n_0_1_26));
   INV_X1 i_0_1_53 (.A(n_0_1_27), .ZN(n_0_60));
   AOI222_X1 i_0_1_54 (.A1(n_0_1_44), .A2(A[20]), .B1(SubM[20]), .B2(n_0_1_42), 
      .C1(AddM[20]), .C2(n_0_1_43), .ZN(n_0_1_27));
   INV_X1 i_0_1_55 (.A(n_0_1_28), .ZN(n_0_61));
   AOI222_X1 i_0_1_56 (.A1(n_0_1_44), .A2(A[21]), .B1(SubM[21]), .B2(n_0_1_42), 
      .C1(AddM[21]), .C2(n_0_1_43), .ZN(n_0_1_28));
   INV_X1 i_0_1_57 (.A(n_0_1_29), .ZN(n_0_62));
   AOI222_X1 i_0_1_58 (.A1(n_0_1_44), .A2(A[22]), .B1(SubM[22]), .B2(n_0_1_42), 
      .C1(AddM[22]), .C2(n_0_1_43), .ZN(n_0_1_29));
   INV_X1 i_0_1_59 (.A(n_0_1_30), .ZN(n_0_63));
   AOI222_X1 i_0_1_60 (.A1(n_0_1_44), .A2(A[23]), .B1(SubM[23]), .B2(n_0_1_42), 
      .C1(AddM[23]), .C2(n_0_1_43), .ZN(n_0_1_30));
   INV_X1 i_0_1_61 (.A(n_0_1_31), .ZN(n_0_64));
   AOI222_X1 i_0_1_62 (.A1(n_0_1_44), .A2(A[24]), .B1(SubM[24]), .B2(n_0_1_42), 
      .C1(AddM[24]), .C2(n_0_1_43), .ZN(n_0_1_31));
   INV_X1 i_0_1_63 (.A(n_0_1_32), .ZN(n_0_65));
   AOI222_X1 i_0_1_64 (.A1(n_0_1_44), .A2(A[25]), .B1(SubM[25]), .B2(n_0_1_42), 
      .C1(AddM[25]), .C2(n_0_1_43), .ZN(n_0_1_32));
   INV_X1 i_0_1_65 (.A(n_0_1_33), .ZN(n_0_66));
   AOI222_X1 i_0_1_66 (.A1(n_0_1_44), .A2(A[26]), .B1(SubM[26]), .B2(n_0_1_42), 
      .C1(AddM[26]), .C2(n_0_1_43), .ZN(n_0_1_33));
   INV_X1 i_0_1_67 (.A(n_0_1_34), .ZN(n_0_67));
   AOI222_X1 i_0_1_68 (.A1(n_0_1_44), .A2(A[27]), .B1(SubM[27]), .B2(n_0_1_42), 
      .C1(AddM[27]), .C2(n_0_1_43), .ZN(n_0_1_34));
   INV_X1 i_0_1_69 (.A(n_0_1_35), .ZN(n_0_68));
   AOI222_X1 i_0_1_70 (.A1(n_0_1_44), .A2(A[28]), .B1(SubM[28]), .B2(n_0_1_42), 
      .C1(AddM[28]), .C2(n_0_1_43), .ZN(n_0_1_35));
   INV_X1 i_0_1_71 (.A(n_0_1_36), .ZN(n_0_69));
   AOI222_X1 i_0_1_72 (.A1(n_0_1_44), .A2(A[29]), .B1(SubM[29]), .B2(n_0_1_42), 
      .C1(AddM[29]), .C2(n_0_1_43), .ZN(n_0_1_36));
   INV_X1 i_0_1_73 (.A(n_0_1_37), .ZN(n_0_70));
   AOI222_X1 i_0_1_74 (.A1(n_0_1_44), .A2(A[30]), .B1(SubM[30]), .B2(n_0_1_42), 
      .C1(AddM[30]), .C2(n_0_1_43), .ZN(n_0_1_37));
   NAND2_X1 i_0_1_75 (.A1(n_0_1_38), .A2(n_0_1_39), .ZN(n_0_71));
   NAND2_X1 i_0_1_76 (.A1(n_0_1_44), .A2(A[31]), .ZN(n_0_1_38));
   INV_X1 i_0_1_77 (.A(n_0_1_39), .ZN(n_0_72));
   AOI22_X1 i_0_1_78 (.A1(AddM[31]), .A2(n_0_1_43), .B1(n_0_1_42), .B2(SubM[31]), 
      .ZN(n_0_1_39));
   MUX2_X1 i_0_1_79 (.A(l8[1]), .B(read2[0]), .S(start), .Z(n_0_104));
   MUX2_X1 i_0_1_80 (.A(l8[2]), .B(read2[1]), .S(start), .Z(n_0_105));
   MUX2_X1 i_0_1_81 (.A(l8[3]), .B(read2[2]), .S(start), .Z(n_0_106));
   MUX2_X1 i_0_1_82 (.A(l8[4]), .B(read2[3]), .S(start), .Z(n_0_107));
   MUX2_X1 i_0_1_83 (.A(l8[5]), .B(read2[4]), .S(start), .Z(n_0_108));
   MUX2_X1 i_0_1_84 (.A(l8[6]), .B(read2[5]), .S(start), .Z(n_0_109));
   MUX2_X1 i_0_1_85 (.A(l8[7]), .B(read2[6]), .S(start), .Z(n_0_73));
   MUX2_X1 i_0_1_86 (.A(l8[8]), .B(read2[7]), .S(start), .Z(n_0_74));
   MUX2_X1 i_0_1_87 (.A(l8[9]), .B(read2[8]), .S(start), .Z(n_0_75));
   MUX2_X1 i_0_1_88 (.A(l8[10]), .B(read2[9]), .S(start), .Z(n_0_76));
   MUX2_X1 i_0_1_89 (.A(l8[11]), .B(read2[10]), .S(start), .Z(n_0_77));
   MUX2_X1 i_0_1_90 (.A(l8[12]), .B(read2[11]), .S(start), .Z(n_0_78));
   MUX2_X1 i_0_1_91 (.A(l8[13]), .B(read2[12]), .S(start), .Z(n_0_79));
   MUX2_X1 i_0_1_92 (.A(l8[14]), .B(read2[13]), .S(start), .Z(n_0_80));
   MUX2_X1 i_0_1_93 (.A(l8[15]), .B(read2[14]), .S(start), .Z(n_0_81));
   MUX2_X1 i_0_1_94 (.A(l8[16]), .B(read2[15]), .S(start), .Z(n_0_82));
   MUX2_X1 i_0_1_95 (.A(l8[17]), .B(read2[16]), .S(start), .Z(n_0_83));
   MUX2_X1 i_0_1_96 (.A(l8[18]), .B(read2[17]), .S(start), .Z(n_0_84));
   MUX2_X1 i_0_1_97 (.A(l8[19]), .B(read2[18]), .S(start), .Z(n_0_85));
   MUX2_X1 i_0_1_98 (.A(l8[20]), .B(read2[19]), .S(start), .Z(n_0_86));
   MUX2_X1 i_0_1_99 (.A(l8[21]), .B(read2[20]), .S(start), .Z(n_0_87));
   MUX2_X1 i_0_1_100 (.A(l8[22]), .B(read2[21]), .S(start), .Z(n_0_88));
   MUX2_X1 i_0_1_101 (.A(l8[23]), .B(read2[22]), .S(start), .Z(n_0_89));
   MUX2_X1 i_0_1_102 (.A(l8[24]), .B(read2[23]), .S(start), .Z(n_0_90));
   MUX2_X1 i_0_1_103 (.A(l8[25]), .B(read2[24]), .S(start), .Z(n_0_91));
   MUX2_X1 i_0_1_104 (.A(l8[26]), .B(read2[25]), .S(start), .Z(n_0_92));
   MUX2_X1 i_0_1_105 (.A(l8[27]), .B(read2[26]), .S(start), .Z(n_0_93));
   MUX2_X1 i_0_1_106 (.A(l8[28]), .B(read2[27]), .S(start), .Z(n_0_94));
   MUX2_X1 i_0_1_107 (.A(l8[29]), .B(read2[28]), .S(start), .Z(n_0_95));
   MUX2_X1 i_0_1_108 (.A(l8[30]), .B(read2[29]), .S(start), .Z(n_0_96));
   MUX2_X1 i_0_1_109 (.A(l8[31]), .B(read2[30]), .S(start), .Z(n_0_97));
   NAND2_X1 i_0_1_110 (.A1(n_0_1_41), .A2(n_0_1_40), .ZN(n_0_98));
   AOI22_X1 i_0_1_111 (.A1(AddM[0]), .A2(n_0_1_43), .B1(n_0_1_42), .B2(SubM[0]), 
      .ZN(n_0_1_40));
   AOI22_X1 i_0_1_112 (.A1(n_0_1_44), .A2(A[0]), .B1(start), .B2(read2[31]), 
      .ZN(n_0_1_41));
   NOR3_X1 i_0_1_113 (.A1(n_0_1_49), .A2(start), .A3(q0), .ZN(n_0_1_42));
   AND3_X1 i_0_1_114 (.A1(n_0_1_49), .A2(n_0_33), .A3(q0), .ZN(n_0_1_43));
   AOI21_X1 i_0_1_115 (.A(n_0_1_44), .B1(n_0_1_46), .B2(n_0_33), .ZN(n_0_101));
   NOR2_X1 i_0_1_116 (.A1(n_0_1_45), .A2(start), .ZN(n_0_1_44));
   XNOR2_X1 i_0_1_117 (.A(q0), .B(n_0_1_49), .ZN(n_0_1_45));
   NOR2_X1 i_0_1_118 (.A1(n_0_1_49), .A2(start), .ZN(n_0_99));
   NAND2_X1 i_0_1_119 (.A1(n_0_1_46), .A2(n_0_33), .ZN(n_0_100));
   NOR4_X1 i_0_1_120 (.A1(n_0_1_47), .A2(count[2]), .A3(count[3]), .A4(count[4]), 
      .ZN(n_0_1_46));
   NAND2_X1 i_0_1_121 (.A1(count[5]), .A2(n_0_1_48), .ZN(n_0_1_47));
   NOR2_X1 i_0_1_122 (.A1(count[1]), .A2(count[0]), .ZN(n_0_1_48));
   INV_X1 i_0_1_123 (.A(start), .ZN(n_0_33));
   INV_X1 i_0_1_124 (.A(l8[0]), .ZN(n_0_1_49));
endmodule
