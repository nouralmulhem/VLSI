/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 13:02:04 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1473625449 */

module subnormal(inputA, inputB, overflow, signal, result);
   input [7:0]inputA;
   input [7:0]inputB;
   output overflow;
   output signal;
   output [31:0]result;

   wire n_32_0_0;
   wire n_32_0_1;
   wire n_32_0_2;
   wire n_32_0_3;
   wire n_32_0_4;
   wire n_32_0_5;
   wire n_32_0_6;
   wire n_32_0_7;
   wire n_32_0_8;

   TBUF_X1 i_0 (.A(1'b0), .EN(n_0), .Z(result[0]));
   TBUF_X1 i_1 (.A(1'b0), .EN(n_0), .Z(result[1]));
   TBUF_X1 i_2 (.A(1'b0), .EN(n_0), .Z(result[2]));
   TBUF_X1 i_3 (.A(1'b0), .EN(n_0), .Z(result[3]));
   TBUF_X1 i_4 (.A(1'b0), .EN(n_0), .Z(result[4]));
   TBUF_X1 i_5 (.A(1'b0), .EN(n_0), .Z(result[5]));
   TBUF_X1 i_6 (.A(1'b0), .EN(n_0), .Z(result[6]));
   TBUF_X1 i_7 (.A(1'b0), .EN(n_0), .Z(result[7]));
   TBUF_X1 i_8 (.A(1'b0), .EN(n_0), .Z(result[8]));
   TBUF_X1 i_9 (.A(1'b0), .EN(n_0), .Z(result[9]));
   TBUF_X1 i_10 (.A(1'b0), .EN(n_0), .Z(result[10]));
   TBUF_X1 i_11 (.A(1'b0), .EN(n_0), .Z(result[11]));
   TBUF_X1 i_12 (.A(1'b0), .EN(n_0), .Z(result[12]));
   TBUF_X1 i_13 (.A(1'b0), .EN(n_0), .Z(result[13]));
   TBUF_X1 i_14 (.A(1'b0), .EN(n_0), .Z(result[14]));
   TBUF_X1 i_15 (.A(1'b0), .EN(n_0), .Z(result[15]));
   TBUF_X1 i_16 (.A(1'b0), .EN(n_0), .Z(result[16]));
   TBUF_X1 i_17 (.A(1'b0), .EN(n_0), .Z(result[17]));
   TBUF_X1 i_18 (.A(1'b0), .EN(n_0), .Z(result[18]));
   TBUF_X1 i_19 (.A(1'b0), .EN(n_0), .Z(result[19]));
   TBUF_X1 i_20 (.A(1'b0), .EN(n_0), .Z(result[20]));
   TBUF_X1 i_21 (.A(1'b0), .EN(n_0), .Z(result[21]));
   TBUF_X1 i_22 (.A(1'b0), .EN(n_0), .Z(result[22]));
   TBUF_X1 i_23 (.A(1'b0), .EN(n_0), .Z(result[23]));
   TBUF_X1 i_24 (.A(1'b0), .EN(n_0), .Z(result[24]));
   TBUF_X1 i_25 (.A(1'b0), .EN(n_0), .Z(result[25]));
   TBUF_X1 i_26 (.A(1'b0), .EN(n_0), .Z(result[26]));
   TBUF_X1 i_27 (.A(1'b0), .EN(n_0), .Z(result[27]));
   TBUF_X1 i_28 (.A(1'b0), .EN(n_0), .Z(result[28]));
   TBUF_X1 i_29 (.A(1'b0), .EN(n_0), .Z(result[29]));
   TBUF_X1 i_30 (.A(1'b0), .EN(n_0), .Z(result[30]));
   TBUF_X1 i_31 (.A(1'b0), .EN(n_0), .Z(result[31]));
   INV_X1 i_32_0_0 (.A(n_32_0_0), .ZN(overflow));
   AOI221_X1 i_32_0_1 (.A(n_0), .B1(n_32_0_4), .B2(n_32_0_3), .C1(n_32_0_2), 
      .C2(n_32_0_1), .ZN(n_32_0_0));
   NOR4_X1 i_32_0_2 (.A1(inputB[7]), .A2(inputB[6]), .A3(inputB[5]), .A4(
      inputB[4]), .ZN(n_32_0_1));
   NOR4_X1 i_32_0_3 (.A1(inputB[3]), .A2(inputB[2]), .A3(inputB[1]), .A4(
      inputB[0]), .ZN(n_32_0_2));
   NOR4_X1 i_32_0_4 (.A1(inputA[7]), .A2(inputA[6]), .A3(inputA[5]), .A4(
      inputA[4]), .ZN(n_32_0_3));
   NOR4_X1 i_32_0_5 (.A1(inputA[3]), .A2(inputA[2]), .A3(inputA[1]), .A4(
      inputA[0]), .ZN(n_32_0_4));
   OAI22_X1 i_32_0_6 (.A1(n_32_0_8), .A2(n_32_0_7), .B1(n_32_0_6), .B2(n_32_0_5), 
      .ZN(n_0));
   NAND4_X1 i_32_0_7 (.A1(inputB[7]), .A2(inputB[6]), .A3(inputB[5]), .A4(
      inputB[4]), .ZN(n_32_0_5));
   NAND4_X1 i_32_0_8 (.A1(inputB[3]), .A2(inputB[2]), .A3(inputB[1]), .A4(
      inputB[0]), .ZN(n_32_0_6));
   NAND4_X1 i_32_0_9 (.A1(inputA[7]), .A2(inputA[6]), .A3(inputA[5]), .A4(
      inputA[4]), .ZN(n_32_0_7));
   NAND4_X1 i_32_0_10 (.A1(inputA[3]), .A2(inputA[2]), .A3(inputA[1]), .A4(
      inputA[0]), .ZN(n_32_0_8));
endmodule

module xor_module(sign1, sign2, sign_out);
   input sign1;
   input sign2;
   output sign_out;

   XOR2_X1 i_0_0 (.A(sign1), .B(sign2), .Z(sign_out));
endmodule

module full_adder__0_88(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
   AND2_X1 i_0_1 (.A1(i_bit2), .A2(i_bit1), .ZN(o_carry));
endmodule

module full_adder__0_84(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_80(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_76(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_72(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_68(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_64(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_60(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module ripple_adder__0_89(i_add1, i_add2, o_result, o_carry);
   input [7:0]i_add1;
   input [7:0]i_add2;
   output [7:0]o_result;
   output o_carry;

   full_adder__0_88 genblk1_0_full_adder_inst (.i_bit1(i_add1[0]), .i_bit2(
      i_add2[0]), .i_carry(), .o_sum(o_result[0]), .o_carry(n_0));
   full_adder__0_84 genblk1_1_full_adder_inst (.i_bit1(i_add1[1]), .i_bit2(
      i_add2[1]), .i_carry(n_0), .o_sum(o_result[1]), .o_carry(n_1));
   full_adder__0_80 genblk1_2_full_adder_inst (.i_bit1(i_add1[2]), .i_bit2(
      i_add2[2]), .i_carry(n_1), .o_sum(o_result[2]), .o_carry(n_2));
   full_adder__0_76 genblk1_3_full_adder_inst (.i_bit1(i_add1[3]), .i_bit2(
      i_add2[3]), .i_carry(n_2), .o_sum(o_result[3]), .o_carry(n_3));
   full_adder__0_72 genblk1_4_full_adder_inst (.i_bit1(i_add1[4]), .i_bit2(
      i_add2[4]), .i_carry(n_3), .o_sum(o_result[4]), .o_carry(n_4));
   full_adder__0_68 genblk1_5_full_adder_inst (.i_bit1(i_add1[5]), .i_bit2(
      i_add2[5]), .i_carry(n_4), .o_sum(o_result[5]), .o_carry(n_5));
   full_adder__0_64 genblk1_6_full_adder_inst (.i_bit1(i_add1[6]), .i_bit2(
      i_add2[6]), .i_carry(n_5), .o_sum(o_result[6]), .o_carry(n_6));
   full_adder__0_60 genblk1_7_full_adder_inst (.i_bit1(i_add1[7]), .i_bit2(
      i_add2[7]), .i_carry(n_6), .o_sum(o_result[7]), .o_carry());
endmodule

module full_adder__0_121(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
   AND2_X1 i_0_1 (.A1(i_bit2), .A2(i_bit1), .ZN(o_carry));
endmodule

module full_adder__0_117(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_113(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_109(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_105(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_101(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_97(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_93(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module ripple_adder__0_122(i_add1, i_add2, o_result, o_carry);
   input [7:0]i_add1;
   input [7:0]i_add2;
   output [7:0]o_result;
   output o_carry;

   full_adder__0_121 genblk1_0_full_adder_inst (.i_bit1(i_add1[0]), .i_bit2(
      i_add2[0]), .i_carry(), .o_sum(o_result[0]), .o_carry(n_0));
   full_adder__0_117 genblk1_1_full_adder_inst (.i_bit1(i_add1[1]), .i_bit2(
      i_add2[1]), .i_carry(n_0), .o_sum(o_result[1]), .o_carry(n_1));
   full_adder__0_113 genblk1_2_full_adder_inst (.i_bit1(i_add1[2]), .i_bit2(
      i_add2[2]), .i_carry(n_1), .o_sum(o_result[2]), .o_carry(n_2));
   full_adder__0_109 genblk1_3_full_adder_inst (.i_bit1(i_add1[3]), .i_bit2(
      i_add2[3]), .i_carry(n_2), .o_sum(o_result[3]), .o_carry(n_3));
   full_adder__0_105 genblk1_4_full_adder_inst (.i_bit1(i_add1[4]), .i_bit2(
      i_add2[4]), .i_carry(n_3), .o_sum(o_result[4]), .o_carry(n_4));
   full_adder__0_101 genblk1_5_full_adder_inst (.i_bit1(i_add1[5]), .i_bit2(
      i_add2[5]), .i_carry(n_4), .o_sum(o_result[5]), .o_carry(n_5));
   full_adder__0_97 genblk1_6_full_adder_inst (.i_bit1(i_add1[6]), .i_bit2(
      i_add2[6]), .i_carry(n_5), .o_sum(o_result[6]), .o_carry(n_6));
   full_adder__0_93 genblk1_7_full_adder_inst (.i_bit1(i_add1[7]), .i_bit2(
      i_add2[7]), .i_carry(n_6), .o_sum(o_result[7]), .o_carry(o_carry));
endmodule

module regFile__0_123(read_data, read_data2, write_en, write_data, write_data2, 
      clk);
   output [24:0]read_data;
   output [24:0]read_data2;
   input write_en;
   input [24:0]write_data;
   input [24:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[22]  (.D(write_data2[22]), .CK(n_0), .Q(read_data2[22]), 
      .QN());
   DFF_X1 \my_reg2_reg[21]  (.D(write_data2[21]), .CK(n_0), .Q(read_data2[21]), 
      .QN());
   DFF_X1 \my_reg2_reg[20]  (.D(write_data2[20]), .CK(n_0), .Q(read_data2[20]), 
      .QN());
   DFF_X1 \my_reg2_reg[19]  (.D(write_data2[19]), .CK(n_0), .Q(read_data2[19]), 
      .QN());
   DFF_X1 \my_reg2_reg[18]  (.D(write_data2[18]), .CK(n_0), .Q(read_data2[18]), 
      .QN());
   DFF_X1 \my_reg2_reg[17]  (.D(write_data2[17]), .CK(n_0), .Q(read_data2[17]), 
      .QN());
   DFF_X1 \my_reg2_reg[16]  (.D(write_data2[16]), .CK(n_0), .Q(read_data2[16]), 
      .QN());
   DFF_X1 \my_reg2_reg[15]  (.D(write_data2[15]), .CK(n_0), .Q(read_data2[15]), 
      .QN());
   DFF_X1 \my_reg2_reg[14]  (.D(write_data2[14]), .CK(n_0), .Q(read_data2[14]), 
      .QN());
   DFF_X1 \my_reg2_reg[13]  (.D(write_data2[13]), .CK(n_0), .Q(read_data2[13]), 
      .QN());
   DFF_X1 \my_reg2_reg[12]  (.D(write_data2[12]), .CK(n_0), .Q(read_data2[12]), 
      .QN());
   DFF_X1 \my_reg2_reg[11]  (.D(write_data2[11]), .CK(n_0), .Q(read_data2[11]), 
      .QN());
   DFF_X1 \my_reg2_reg[10]  (.D(write_data2[10]), .CK(n_0), .Q(read_data2[10]), 
      .QN());
   DFF_X1 \my_reg2_reg[9]  (.D(write_data2[9]), .CK(n_0), .Q(read_data2[9]), 
      .QN());
   DFF_X1 \my_reg2_reg[8]  (.D(write_data2[8]), .CK(n_0), .Q(read_data2[8]), 
      .QN());
   DFF_X1 \my_reg2_reg[7]  (.D(write_data2[7]), .CK(n_0), .Q(read_data2[7]), 
      .QN());
   DFF_X1 \my_reg2_reg[6]  (.D(write_data2[6]), .CK(n_0), .Q(read_data2[6]), 
      .QN());
   DFF_X1 \my_reg2_reg[5]  (.D(write_data2[5]), .CK(n_0), .Q(read_data2[5]), 
      .QN());
   DFF_X1 \my_reg2_reg[4]  (.D(write_data2[4]), .CK(n_0), .Q(read_data2[4]), 
      .QN());
   DFF_X1 \my_reg2_reg[3]  (.D(write_data2[3]), .CK(n_0), .Q(read_data2[3]), 
      .QN());
   DFF_X1 \my_reg2_reg[2]  (.D(write_data2[2]), .CK(n_0), .Q(read_data2[2]), 
      .QN());
   DFF_X1 \my_reg2_reg[1]  (.D(write_data2[1]), .CK(n_0), .Q(read_data2[1]), 
      .QN());
   DFF_X1 \my_reg2_reg[0]  (.D(write_data2[0]), .CK(n_0), .Q(read_data2[0]), 
      .QN());
   DFF_X1 \my_reg_reg[22]  (.D(write_data[22]), .CK(n_0), .Q(read_data[22]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg2_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
   DFF_X1 \my_reg2_reg[24]  (.D(write_data[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
endmodule

module fullAdder__0_420(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_414(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_411(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_408(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_405(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_402(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_399(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_396(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_393(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_390(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_387(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_384(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_381(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_378(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_375(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_372(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_369(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_366(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_363(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_360(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_357(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_354(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_351(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_348(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_345(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_342(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(y), .B(x), .Z(sum));
endmodule

module fullAdder__0_339(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_336(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_333(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_330(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_327(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_324(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_321(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_318(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_315(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_312(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_309(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_306(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_303(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_300(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_297(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_294(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_291(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_288(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_285(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_282(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_279(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_276(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_273(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(x), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(y), .ZN(sum));
endmodule

module carrySaveAdder__0_421(a, b, c, sum, cout);
   input [24:0]a;
   input [24:0]b;
   input [24:0]c;
   output [24:0]sum;
   output cout;

   wire [24:0]halfcarry;
   wire [24:0]halfcout;
   wire [24:0]halfsum;

   fullAdder__0_420 fulladder_f2 (.x(halfsum[1]), .y(halfcout[0]), .cin(), 
      .sum(sum[1]), .cout(halfcarry[0]));
   fullAdder__0_414 genblk1_0_fulladder_f1 (.x(a[0]), .y(b[0]), .cin(), .sum(
      sum[0]), .cout(halfcout[0]));
   fullAdder__0_411 genblk1_1_fulladder_f1 (.x(a[1]), .y(b[1]), .cin(), .sum(
      halfsum[1]), .cout(halfcout[1]));
   fullAdder__0_408 genblk1_2_fulladder_f1 (.x(a[2]), .y(b[2]), .cin(), .sum(
      halfsum[2]), .cout(halfcout[2]));
   fullAdder__0_405 genblk1_3_fulladder_f1 (.x(a[3]), .y(b[3]), .cin(), .sum(
      halfsum[3]), .cout(halfcout[3]));
   fullAdder__0_402 genblk1_4_fulladder_f1 (.x(a[4]), .y(b[4]), .cin(), .sum(
      halfsum[4]), .cout(halfcout[4]));
   fullAdder__0_399 genblk1_5_fulladder_f1 (.x(a[5]), .y(b[5]), .cin(), .sum(
      halfsum[5]), .cout(halfcout[5]));
   fullAdder__0_396 genblk1_6_fulladder_f1 (.x(a[6]), .y(b[6]), .cin(), .sum(
      halfsum[6]), .cout(halfcout[6]));
   fullAdder__0_393 genblk1_7_fulladder_f1 (.x(a[7]), .y(b[7]), .cin(), .sum(
      halfsum[7]), .cout(halfcout[7]));
   fullAdder__0_390 genblk1_8_fulladder_f1 (.x(a[8]), .y(b[8]), .cin(), .sum(
      halfsum[8]), .cout(halfcout[8]));
   fullAdder__0_387 genblk1_9_fulladder_f1 (.x(a[9]), .y(b[9]), .cin(), .sum(
      halfsum[9]), .cout(halfcout[9]));
   fullAdder__0_384 genblk1_10_fulladder_f1 (.x(a[10]), .y(b[10]), .cin(), 
      .sum(halfsum[10]), .cout(halfcout[10]));
   fullAdder__0_381 genblk1_11_fulladder_f1 (.x(a[11]), .y(b[11]), .cin(), 
      .sum(halfsum[11]), .cout(halfcout[11]));
   fullAdder__0_378 genblk1_12_fulladder_f1 (.x(a[12]), .y(b[12]), .cin(), 
      .sum(halfsum[12]), .cout(halfcout[12]));
   fullAdder__0_375 genblk1_13_fulladder_f1 (.x(a[13]), .y(b[13]), .cin(), 
      .sum(halfsum[13]), .cout(halfcout[13]));
   fullAdder__0_372 genblk1_14_fulladder_f1 (.x(a[14]), .y(b[14]), .cin(), 
      .sum(halfsum[14]), .cout(halfcout[14]));
   fullAdder__0_369 genblk1_15_fulladder_f1 (.x(a[15]), .y(b[15]), .cin(), 
      .sum(halfsum[15]), .cout(halfcout[15]));
   fullAdder__0_366 genblk1_16_fulladder_f1 (.x(a[16]), .y(b[16]), .cin(), 
      .sum(halfsum[16]), .cout(halfcout[16]));
   fullAdder__0_363 genblk1_17_fulladder_f1 (.x(a[17]), .y(b[17]), .cin(), 
      .sum(halfsum[17]), .cout(halfcout[17]));
   fullAdder__0_360 genblk1_18_fulladder_f1 (.x(a[18]), .y(b[18]), .cin(), 
      .sum(halfsum[18]), .cout(halfcout[18]));
   fullAdder__0_357 genblk1_19_fulladder_f1 (.x(a[19]), .y(b[19]), .cin(), 
      .sum(halfsum[19]), .cout(halfcout[19]));
   fullAdder__0_354 genblk1_20_fulladder_f1 (.x(a[20]), .y(b[20]), .cin(), 
      .sum(halfsum[20]), .cout(halfcout[20]));
   fullAdder__0_351 genblk1_21_fulladder_f1 (.x(a[21]), .y(b[21]), .cin(), 
      .sum(halfsum[21]), .cout(halfcout[21]));
   fullAdder__0_348 genblk1_22_fulladder_f1 (.x(a[22]), .y(b[22]), .cin(), 
      .sum(halfsum[22]), .cout(halfcout[22]));
   fullAdder__0_345 genblk1_23_fulladder_f1 (.x(a[23]), .y(b[23]), .cin(), 
      .sum(halfsum[23]), .cout(halfcout[23]));
   fullAdder__0_342 genblk1_24_fulladder_f1 (.x(a[24]), .y(b[24]), .cin(), 
      .sum(halfsum[24]), .cout());
   fullAdder__0_339 genblk2_1_f3 (.x(halfsum[2]), .y(halfcout[1]), .cin(
      halfcarry[0]), .sum(sum[2]), .cout(halfcarry[1]));
   fullAdder__0_336 genblk2_2_f3 (.x(halfsum[3]), .y(halfcout[2]), .cin(
      halfcarry[1]), .sum(sum[3]), .cout(halfcarry[2]));
   fullAdder__0_333 genblk2_3_f3 (.x(halfsum[4]), .y(halfcout[3]), .cin(
      halfcarry[2]), .sum(sum[4]), .cout(halfcarry[3]));
   fullAdder__0_330 genblk2_4_f3 (.x(halfsum[5]), .y(halfcout[4]), .cin(
      halfcarry[3]), .sum(sum[5]), .cout(halfcarry[4]));
   fullAdder__0_327 genblk2_5_f3 (.x(halfsum[6]), .y(halfcout[5]), .cin(
      halfcarry[4]), .sum(sum[6]), .cout(halfcarry[5]));
   fullAdder__0_324 genblk2_6_f3 (.x(halfsum[7]), .y(halfcout[6]), .cin(
      halfcarry[5]), .sum(sum[7]), .cout(halfcarry[6]));
   fullAdder__0_321 genblk2_7_f3 (.x(halfsum[8]), .y(halfcout[7]), .cin(
      halfcarry[6]), .sum(sum[8]), .cout(halfcarry[7]));
   fullAdder__0_318 genblk2_8_f3 (.x(halfsum[9]), .y(halfcout[8]), .cin(
      halfcarry[7]), .sum(sum[9]), .cout(halfcarry[8]));
   fullAdder__0_315 genblk2_9_f3 (.x(halfsum[10]), .y(halfcout[9]), .cin(
      halfcarry[8]), .sum(sum[10]), .cout(halfcarry[9]));
   fullAdder__0_312 genblk2_10_f3 (.x(halfsum[11]), .y(halfcout[10]), .cin(
      halfcarry[9]), .sum(sum[11]), .cout(halfcarry[10]));
   fullAdder__0_309 genblk2_11_f3 (.x(halfsum[12]), .y(halfcout[11]), .cin(
      halfcarry[10]), .sum(sum[12]), .cout(halfcarry[11]));
   fullAdder__0_306 genblk2_12_f3 (.x(halfsum[13]), .y(halfcout[12]), .cin(
      halfcarry[11]), .sum(sum[13]), .cout(halfcarry[12]));
   fullAdder__0_303 genblk2_13_f3 (.x(halfsum[14]), .y(halfcout[13]), .cin(
      halfcarry[12]), .sum(sum[14]), .cout(halfcarry[13]));
   fullAdder__0_300 genblk2_14_f3 (.x(halfsum[15]), .y(halfcout[14]), .cin(
      halfcarry[13]), .sum(sum[15]), .cout(halfcarry[14]));
   fullAdder__0_297 genblk2_15_f3 (.x(halfsum[16]), .y(halfcout[15]), .cin(
      halfcarry[14]), .sum(sum[16]), .cout(halfcarry[15]));
   fullAdder__0_294 genblk2_16_f3 (.x(halfsum[17]), .y(halfcout[16]), .cin(
      halfcarry[15]), .sum(sum[17]), .cout(halfcarry[16]));
   fullAdder__0_291 genblk2_17_f3 (.x(halfsum[18]), .y(halfcout[17]), .cin(
      halfcarry[16]), .sum(sum[18]), .cout(halfcarry[17]));
   fullAdder__0_288 genblk2_18_f3 (.x(halfsum[19]), .y(halfcout[18]), .cin(
      halfcarry[17]), .sum(sum[19]), .cout(halfcarry[18]));
   fullAdder__0_285 genblk2_19_f3 (.x(halfsum[20]), .y(halfcout[19]), .cin(
      halfcarry[18]), .sum(sum[20]), .cout(halfcarry[19]));
   fullAdder__0_282 genblk2_20_f3 (.x(halfsum[21]), .y(halfcout[20]), .cin(
      halfcarry[19]), .sum(sum[21]), .cout(halfcarry[20]));
   fullAdder__0_279 genblk2_21_f3 (.x(halfsum[22]), .y(halfcout[21]), .cin(
      halfcarry[20]), .sum(sum[22]), .cout(halfcarry[21]));
   fullAdder__0_276 genblk2_22_f3 (.x(halfsum[23]), .y(halfcout[22]), .cin(
      halfcarry[21]), .sum(sum[23]), .cout(halfcarry[22]));
   fullAdder__0_273 genblk2_23_f3 (.x(halfsum[24]), .y(halfcout[23]), .cin(
      halfcarry[22]), .sum(sum[24]), .cout());
endmodule

module fullAdder__0_126(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_132(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_135(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_138(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_141(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_144(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_147(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_150(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_153(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_156(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_159(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_162(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_165(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_168(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_171(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_174(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_177(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_180(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_183(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_186(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_189(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_192(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_195(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_198(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_201(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(x), .B(y), .Z(sum));
   AND2_X1 i_0_1 (.A1(y), .A2(x), .ZN(cout));
endmodule

module fullAdder__0_204(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(y), .B(x), .Z(sum));
endmodule

module fullAdder__0_207(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_210(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_213(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_216(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_219(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_222(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_225(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_228(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_231(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_234(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_237(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_240(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_243(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_246(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_249(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_252(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_255(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_258(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_261(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_264(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_267(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder__0_270(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(cout));
   OAI21_X1 i_0_1 (.A(y), .B1(cin), .B2(x), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(y), .B(n_0_1), .ZN(sum));
   XNOR2_X1 i_0_3 (.A(cin), .B(x), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(cin), .A2(x), .ZN(n_0_2));
endmodule

module fullAdder(x, y, cin, sum, cout);
   input x;
   input y;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(x), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(n_0_0), .B(y), .ZN(sum));
endmodule

module carrySaveAdder(a, b, c, sum, cout);
   input [24:0]a;
   input [24:0]b;
   input [24:0]c;
   output [24:0]sum;
   output cout;

   wire [24:0]halfcarry;
   wire [24:0]halfcout;
   wire [24:0]halfsum;

   fullAdder__0_126 fulladder_f2 (.x(halfsum[1]), .y(halfcout[0]), .cin(), 
      .sum(sum[1]), .cout(halfcarry[0]));
   fullAdder__0_132 genblk1_0_fulladder_f1 (.x(a[0]), .y(b[0]), .cin(), .sum(
      sum[0]), .cout(halfcout[0]));
   fullAdder__0_135 genblk1_1_fulladder_f1 (.x(a[1]), .y(b[1]), .cin(), .sum(
      halfsum[1]), .cout(halfcout[1]));
   fullAdder__0_138 genblk1_2_fulladder_f1 (.x(a[2]), .y(b[2]), .cin(), .sum(
      halfsum[2]), .cout(halfcout[2]));
   fullAdder__0_141 genblk1_3_fulladder_f1 (.x(a[3]), .y(b[3]), .cin(), .sum(
      halfsum[3]), .cout(halfcout[3]));
   fullAdder__0_144 genblk1_4_fulladder_f1 (.x(a[4]), .y(b[4]), .cin(), .sum(
      halfsum[4]), .cout(halfcout[4]));
   fullAdder__0_147 genblk1_5_fulladder_f1 (.x(a[5]), .y(b[5]), .cin(), .sum(
      halfsum[5]), .cout(halfcout[5]));
   fullAdder__0_150 genblk1_6_fulladder_f1 (.x(a[6]), .y(b[6]), .cin(), .sum(
      halfsum[6]), .cout(halfcout[6]));
   fullAdder__0_153 genblk1_7_fulladder_f1 (.x(a[7]), .y(b[7]), .cin(), .sum(
      halfsum[7]), .cout(halfcout[7]));
   fullAdder__0_156 genblk1_8_fulladder_f1 (.x(a[8]), .y(b[8]), .cin(), .sum(
      halfsum[8]), .cout(halfcout[8]));
   fullAdder__0_159 genblk1_9_fulladder_f1 (.x(a[9]), .y(b[9]), .cin(), .sum(
      halfsum[9]), .cout(halfcout[9]));
   fullAdder__0_162 genblk1_10_fulladder_f1 (.x(a[10]), .y(b[10]), .cin(), 
      .sum(halfsum[10]), .cout(halfcout[10]));
   fullAdder__0_165 genblk1_11_fulladder_f1 (.x(a[11]), .y(b[11]), .cin(), 
      .sum(halfsum[11]), .cout(halfcout[11]));
   fullAdder__0_168 genblk1_12_fulladder_f1 (.x(a[12]), .y(b[12]), .cin(), 
      .sum(halfsum[12]), .cout(halfcout[12]));
   fullAdder__0_171 genblk1_13_fulladder_f1 (.x(a[13]), .y(b[13]), .cin(), 
      .sum(halfsum[13]), .cout(halfcout[13]));
   fullAdder__0_174 genblk1_14_fulladder_f1 (.x(a[14]), .y(b[14]), .cin(), 
      .sum(halfsum[14]), .cout(halfcout[14]));
   fullAdder__0_177 genblk1_15_fulladder_f1 (.x(a[15]), .y(b[15]), .cin(), 
      .sum(halfsum[15]), .cout(halfcout[15]));
   fullAdder__0_180 genblk1_16_fulladder_f1 (.x(a[16]), .y(b[16]), .cin(), 
      .sum(halfsum[16]), .cout(halfcout[16]));
   fullAdder__0_183 genblk1_17_fulladder_f1 (.x(a[17]), .y(b[17]), .cin(), 
      .sum(halfsum[17]), .cout(halfcout[17]));
   fullAdder__0_186 genblk1_18_fulladder_f1 (.x(a[18]), .y(b[18]), .cin(), 
      .sum(halfsum[18]), .cout(halfcout[18]));
   fullAdder__0_189 genblk1_19_fulladder_f1 (.x(a[19]), .y(b[19]), .cin(), 
      .sum(halfsum[19]), .cout(halfcout[19]));
   fullAdder__0_192 genblk1_20_fulladder_f1 (.x(a[20]), .y(b[20]), .cin(), 
      .sum(halfsum[20]), .cout(halfcout[20]));
   fullAdder__0_195 genblk1_21_fulladder_f1 (.x(a[21]), .y(b[21]), .cin(), 
      .sum(halfsum[21]), .cout(halfcout[21]));
   fullAdder__0_198 genblk1_22_fulladder_f1 (.x(a[22]), .y(b[22]), .cin(), 
      .sum(halfsum[22]), .cout(halfcout[22]));
   fullAdder__0_201 genblk1_23_fulladder_f1 (.x(a[23]), .y(b[23]), .cin(), 
      .sum(halfsum[23]), .cout(halfcout[23]));
   fullAdder__0_204 genblk1_24_fulladder_f1 (.x(a[24]), .y(b[24]), .cin(), 
      .sum(halfsum[24]), .cout());
   fullAdder__0_207 genblk2_1_f3 (.x(halfsum[2]), .y(halfcout[1]), .cin(
      halfcarry[0]), .sum(sum[2]), .cout(halfcarry[1]));
   fullAdder__0_210 genblk2_2_f3 (.x(halfsum[3]), .y(halfcout[2]), .cin(
      halfcarry[1]), .sum(sum[3]), .cout(halfcarry[2]));
   fullAdder__0_213 genblk2_3_f3 (.x(halfsum[4]), .y(halfcout[3]), .cin(
      halfcarry[2]), .sum(sum[4]), .cout(halfcarry[3]));
   fullAdder__0_216 genblk2_4_f3 (.x(halfsum[5]), .y(halfcout[4]), .cin(
      halfcarry[3]), .sum(sum[5]), .cout(halfcarry[4]));
   fullAdder__0_219 genblk2_5_f3 (.x(halfsum[6]), .y(halfcout[5]), .cin(
      halfcarry[4]), .sum(sum[6]), .cout(halfcarry[5]));
   fullAdder__0_222 genblk2_6_f3 (.x(halfsum[7]), .y(halfcout[6]), .cin(
      halfcarry[5]), .sum(sum[7]), .cout(halfcarry[6]));
   fullAdder__0_225 genblk2_7_f3 (.x(halfsum[8]), .y(halfcout[7]), .cin(
      halfcarry[6]), .sum(sum[8]), .cout(halfcarry[7]));
   fullAdder__0_228 genblk2_8_f3 (.x(halfsum[9]), .y(halfcout[8]), .cin(
      halfcarry[7]), .sum(sum[9]), .cout(halfcarry[8]));
   fullAdder__0_231 genblk2_9_f3 (.x(halfsum[10]), .y(halfcout[9]), .cin(
      halfcarry[8]), .sum(sum[10]), .cout(halfcarry[9]));
   fullAdder__0_234 genblk2_10_f3 (.x(halfsum[11]), .y(halfcout[10]), .cin(
      halfcarry[9]), .sum(sum[11]), .cout(halfcarry[10]));
   fullAdder__0_237 genblk2_11_f3 (.x(halfsum[12]), .y(halfcout[11]), .cin(
      halfcarry[10]), .sum(sum[12]), .cout(halfcarry[11]));
   fullAdder__0_240 genblk2_12_f3 (.x(halfsum[13]), .y(halfcout[12]), .cin(
      halfcarry[11]), .sum(sum[13]), .cout(halfcarry[12]));
   fullAdder__0_243 genblk2_13_f3 (.x(halfsum[14]), .y(halfcout[13]), .cin(
      halfcarry[12]), .sum(sum[14]), .cout(halfcarry[13]));
   fullAdder__0_246 genblk2_14_f3 (.x(halfsum[15]), .y(halfcout[14]), .cin(
      halfcarry[13]), .sum(sum[15]), .cout(halfcarry[14]));
   fullAdder__0_249 genblk2_15_f3 (.x(halfsum[16]), .y(halfcout[15]), .cin(
      halfcarry[14]), .sum(sum[16]), .cout(halfcarry[15]));
   fullAdder__0_252 genblk2_16_f3 (.x(halfsum[17]), .y(halfcout[16]), .cin(
      halfcarry[15]), .sum(sum[17]), .cout(halfcarry[16]));
   fullAdder__0_255 genblk2_17_f3 (.x(halfsum[18]), .y(halfcout[17]), .cin(
      halfcarry[16]), .sum(sum[18]), .cout(halfcarry[17]));
   fullAdder__0_258 genblk2_18_f3 (.x(halfsum[19]), .y(halfcout[18]), .cin(
      halfcarry[17]), .sum(sum[19]), .cout(halfcarry[18]));
   fullAdder__0_261 genblk2_19_f3 (.x(halfsum[20]), .y(halfcout[19]), .cin(
      halfcarry[18]), .sum(sum[20]), .cout(halfcarry[19]));
   fullAdder__0_264 genblk2_20_f3 (.x(halfsum[21]), .y(halfcout[20]), .cin(
      halfcarry[19]), .sum(sum[21]), .cout(halfcarry[20]));
   fullAdder__0_267 genblk2_21_f3 (.x(halfsum[22]), .y(halfcout[21]), .cin(
      halfcarry[20]), .sum(sum[22]), .cout(halfcarry[21]));
   fullAdder__0_270 genblk2_22_f3 (.x(halfsum[23]), .y(halfcout[22]), .cin(
      halfcarry[21]), .sum(sum[23]), .cout(halfcarry[22]));
   fullAdder genblk2_23_f3 (.x(halfsum[24]), .y(halfcout[23]), .cin(
      halfcarry[22]), .sum(sum[24]), .cout());
endmodule

module regFile(read_data, read_data2, write_en, write_data, write_data2, clk);
   output [24:0]read_data;
   output [24:0]read_data2;
   input write_en;
   input [24:0]write_data;
   input [24:0]write_data2;
   input clk;

   DFF_X1 \my_reg2_reg[24]  (.D(write_data2[24]), .CK(n_0), .Q(read_data2[24]), 
      .QN());
   DFF_X1 \my_reg2_reg[23]  (.D(write_data2[23]), .CK(n_0), .Q(read_data2[23]), 
      .QN());
   DFF_X1 \my_reg_reg[21]  (.D(write_data[21]), .CK(n_0), .Q(read_data[21]), 
      .QN());
   DFF_X1 \my_reg_reg[20]  (.D(write_data[20]), .CK(n_0), .Q(read_data[20]), 
      .QN());
   DFF_X1 \my_reg_reg[19]  (.D(write_data[19]), .CK(n_0), .Q(read_data[19]), 
      .QN());
   DFF_X1 \my_reg_reg[18]  (.D(write_data[18]), .CK(n_0), .Q(read_data[18]), 
      .QN());
   DFF_X1 \my_reg_reg[17]  (.D(write_data[17]), .CK(n_0), .Q(read_data[17]), 
      .QN());
   DFF_X1 \my_reg_reg[16]  (.D(write_data[16]), .CK(n_0), .Q(read_data[16]), 
      .QN());
   DFF_X1 \my_reg_reg[15]  (.D(write_data[15]), .CK(n_0), .Q(read_data[15]), 
      .QN());
   DFF_X1 \my_reg_reg[14]  (.D(write_data[14]), .CK(n_0), .Q(read_data[14]), 
      .QN());
   DFF_X1 \my_reg_reg[13]  (.D(write_data[13]), .CK(n_0), .Q(read_data[13]), 
      .QN());
   DFF_X1 \my_reg_reg[12]  (.D(write_data[12]), .CK(n_0), .Q(read_data[12]), 
      .QN());
   DFF_X1 \my_reg_reg[11]  (.D(write_data[11]), .CK(n_0), .Q(read_data[11]), 
      .QN());
   DFF_X1 \my_reg_reg[10]  (.D(write_data[10]), .CK(n_0), .Q(read_data[10]), 
      .QN());
   DFF_X1 \my_reg_reg[9]  (.D(write_data[9]), .CK(n_0), .Q(read_data[9]), .QN());
   DFF_X1 \my_reg_reg[8]  (.D(write_data[8]), .CK(n_0), .Q(read_data[8]), .QN());
   DFF_X1 \my_reg_reg[7]  (.D(write_data[7]), .CK(n_0), .Q(read_data[7]), .QN());
   DFF_X1 \my_reg_reg[6]  (.D(write_data[6]), .CK(n_0), .Q(read_data[6]), .QN());
   DFF_X1 \my_reg_reg[5]  (.D(write_data[5]), .CK(n_0), .Q(read_data[5]), .QN());
   DFF_X1 \my_reg_reg[4]  (.D(write_data[4]), .CK(n_0), .Q(read_data[4]), .QN());
   DFF_X1 \my_reg_reg[3]  (.D(write_data[3]), .CK(n_0), .Q(read_data[3]), .QN());
   DFF_X1 \my_reg_reg[2]  (.D(write_data[2]), .CK(n_0), .Q(read_data[2]), .QN());
   DFF_X1 \my_reg_reg[1]  (.D(write_data[1]), .CK(n_0), .Q(read_data[1]), .QN());
   DFF_X1 \my_reg_reg[0]  (.D(write_data[0]), .CK(n_0), .Q(read_data[0]), .QN());
   CLKGATETST_X1 clk_gate_my_reg_reg (.CK(clk), .E(write_en), .SE(1'b0), 
      .GCK(n_0));
endmodule

module datapath__0_24(f8, p_0);
   input [24:0]f8;
   output [24:0]p_0;

   XOR2_X1 i_0 (.A(f8[1]), .B(f8[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_22), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(f8[2]), .B1(f8[1]), .B2(f8[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(f8[3]), .B(n_22), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(f8[4]), .B(n_21), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(f8[5]), .B(n_20), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_19), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(f8[6]), .B1(n_20), .B2(f8[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(f8[7]), .B(n_19), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(f8[8]), .B(n_18), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_17), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(f8[9]), .B1(n_18), .B2(f8[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(f8[10]), .B(n_17), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(f8[11]), .B(n_16), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(f8[12]), .B(n_15), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(f8[13]), .B(n_14), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(f8[14]), .B(n_13), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(f8[15]), .B(n_12), .Z(p_0[15]));
   XNOR2_X1 i_18 (.A(f8[16]), .B(n_11), .ZN(p_0[16]));
   XOR2_X1 i_19 (.A(f8[17]), .B(n_10), .Z(p_0[17]));
   XOR2_X1 i_20 (.A(f8[18]), .B(n_9), .Z(p_0[18]));
   XOR2_X1 i_21 (.A(f8[19]), .B(n_8), .Z(p_0[19]));
   XNOR2_X1 i_22 (.A(f8[20]), .B(n_7), .ZN(p_0[20]));
   XNOR2_X1 i_23 (.A(f8[21]), .B(n_6), .ZN(p_0[21]));
   XOR2_X1 i_24 (.A(f8[22]), .B(n_5), .Z(p_0[22]));
   XNOR2_X1 i_25 (.A(f8[23]), .B(n_4), .ZN(p_0[23]));
   XNOR2_X1 i_26 (.A(f8[24]), .B(n_3), .ZN(p_0[24]));
   NOR3_X1 i_27 (.A1(n_5), .A2(f8[22]), .A3(f8[23]), .ZN(n_3));
   NOR2_X1 i_28 (.A1(n_5), .A2(f8[22]), .ZN(n_4));
   NAND2_X1 i_29 (.A1(n_6), .A2(n_26), .ZN(n_5));
   NOR3_X1 i_30 (.A1(n_8), .A2(f8[19]), .A3(f8[20]), .ZN(n_6));
   NOR2_X1 i_31 (.A1(n_8), .A2(f8[19]), .ZN(n_7));
   OR2_X1 i_32 (.A1(n_9), .A2(f8[18]), .ZN(n_8));
   OR2_X1 i_33 (.A1(n_10), .A2(f8[17]), .ZN(n_9));
   NAND2_X1 i_34 (.A1(n_11), .A2(n_25), .ZN(n_10));
   NOR2_X1 i_35 (.A1(n_12), .A2(f8[15]), .ZN(n_11));
   NAND2_X1 i_36 (.A1(n_13), .A2(n_24), .ZN(n_12));
   NOR3_X1 i_37 (.A1(n_15), .A2(f8[12]), .A3(f8[13]), .ZN(n_13));
   NOR2_X1 i_38 (.A1(n_15), .A2(f8[12]), .ZN(n_14));
   NAND2_X1 i_39 (.A1(n_16), .A2(n_23), .ZN(n_15));
   NOR2_X1 i_40 (.A1(n_17), .A2(f8[10]), .ZN(n_16));
   OR3_X1 i_41 (.A1(n_18), .A2(f8[8]), .A3(f8[9]), .ZN(n_17));
   OR2_X1 i_42 (.A1(n_19), .A2(f8[7]), .ZN(n_18));
   OR3_X1 i_43 (.A1(n_20), .A2(f8[5]), .A3(f8[6]), .ZN(n_19));
   OR2_X1 i_44 (.A1(n_21), .A2(f8[4]), .ZN(n_20));
   OR2_X1 i_45 (.A1(n_22), .A2(f8[3]), .ZN(n_21));
   OR3_X1 i_46 (.A1(f8[2]), .A2(f8[1]), .A3(f8[0]), .ZN(n_22));
   INV_X1 i_47 (.A(f8[11]), .ZN(n_23));
   INV_X1 i_48 (.A(f8[14]), .ZN(n_24));
   INV_X1 i_49 (.A(f8[16]), .ZN(n_25));
   INV_X1 i_50 (.A(f8[21]), .ZN(n_26));
endmodule

module BoothAlgo(M, Q, result, clk, start);
   input [24:0]M;
   input [24:0]Q;
   output [49:0]result;
   input clk;
   input start;

   wire [24:0]read2;
   wire [24:0]read;
   wire [24:0]SubM;
   wire [24:0]AddM;
   wire [24:0]A;
   wire [24:0]l8;
   wire [24:0]f8;
   wire write_en;
   wire write_en2;
   wire [5:0]count;
   wire q0;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;

   regFile__0_123 inst1 (.read_data({uc_0, uc_1, read[22], read[21], read[20], 
      read[19], read[18], read[17], read[16], read[15], read[14], read[13], 
      read[12], read[11], read[10], read[9], read[8], read[7], read[6], read[5], 
      read[4], read[3], read[2], read[1], read[0]}), .read_data2(read2), 
      .write_en(write_en), .write_data(M), .write_data2({uc_2, uc_3, Q[22], 
      Q[21], Q[20], Q[19], Q[18], Q[17], Q[16], Q[15], Q[14], Q[13], Q[12], 
      Q[11], Q[10], Q[9], Q[8], Q[7], Q[6], Q[5], Q[4], Q[3], Q[2], Q[1], Q[0]}), 
      .clk(clk));
   carrySaveAdder__0_421 subtractor (.a(A), .b({n_86, n_85, n_84, n_58, n_57, 
      n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
      n_44, n_43, n_42, n_41, n_40, n_39, n_38, f8[0]}), .c(), .sum(SubM), .cout());
   carrySaveAdder adder (.a(A), .b(f8), .c(), .sum(AddM), .cout());
   regFile inst2 (.read_data({uc_4, uc_5, uc_6, result[46], result[45], 
      result[44], result[43], result[42], result[41], result[40], result[39], 
      result[38], result[37], result[36], result[35], result[34], result[33], 
      result[32], result[31], result[30], result[29], result[28], result[27], 
      result[26], result[25]}), .read_data2({result[24], result[23], uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29}), 
      .write_en(write_en2), .write_data({uc_30, uc_31, uc_32, A[21], A[20], 
      A[19], A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], A[10], A[9], 
      A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0]}), .write_data2({
      l8[24], l8[23], uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, 
      uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, 
      uc_51, uc_52, uc_53, uc_54, uc_55}), .clk(clk));
   DFF_X1 \A_reg[23]  (.D(n_32), .CK(n_3), .Q(A[23]), .QN());
   DFF_X1 \A_reg[22]  (.D(n_31), .CK(n_3), .Q(A[22]), .QN());
   DFF_X1 \A_reg[21]  (.D(n_30), .CK(n_3), .Q(A[21]), .QN());
   DFF_X1 \A_reg[20]  (.D(n_29), .CK(n_3), .Q(A[20]), .QN());
   DFF_X1 \A_reg[19]  (.D(n_28), .CK(n_3), .Q(A[19]), .QN());
   DFF_X1 \A_reg[18]  (.D(n_27), .CK(n_3), .Q(A[18]), .QN());
   DFF_X1 \A_reg[17]  (.D(n_26), .CK(n_3), .Q(A[17]), .QN());
   DFF_X1 \A_reg[16]  (.D(n_25), .CK(n_3), .Q(A[16]), .QN());
   DFF_X1 \A_reg[15]  (.D(n_24), .CK(n_3), .Q(A[15]), .QN());
   DFF_X1 \A_reg[14]  (.D(n_23), .CK(n_3), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(n_22), .CK(n_3), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(n_21), .CK(n_3), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(n_20), .CK(n_3), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(n_19), .CK(n_3), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(n_18), .CK(n_3), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(n_17), .CK(n_3), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(n_16), .CK(n_3), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(n_15), .CK(n_3), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(n_14), .CK(n_3), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(n_13), .CK(n_3), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(n_12), .CK(n_3), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(n_11), .CK(n_3), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(n_10), .CK(n_3), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(n_9), .CK(n_3), .Q(A[0]), .QN());
   DFF_X1 \A_reg[24]  (.D(n_87), .CK(clk), .Q(A[24]), .QN());
   DFF_X1 \l8_reg[24]  (.D(n_79), .CK(n_3), .Q(l8[24]), .QN());
   DFF_X1 \l8_reg[23]  (.D(n_78), .CK(n_3), .Q(l8[23]), .QN());
   DFF_X1 \l8_reg[22]  (.D(n_77), .CK(n_3), .Q(l8[22]), .QN());
   DFF_X1 \l8_reg[21]  (.D(n_76), .CK(n_3), .Q(l8[21]), .QN());
   DFF_X1 \l8_reg[20]  (.D(n_75), .CK(n_3), .Q(l8[20]), .QN());
   DFF_X1 \l8_reg[19]  (.D(n_74), .CK(n_3), .Q(l8[19]), .QN());
   DFF_X1 \l8_reg[18]  (.D(n_73), .CK(n_3), .Q(l8[18]), .QN());
   DFF_X1 \l8_reg[17]  (.D(n_72), .CK(n_3), .Q(l8[17]), .QN());
   DFF_X1 \l8_reg[16]  (.D(n_71), .CK(n_3), .Q(l8[16]), .QN());
   DFF_X1 \l8_reg[15]  (.D(n_70), .CK(n_3), .Q(l8[15]), .QN());
   DFF_X1 \l8_reg[14]  (.D(n_69), .CK(n_3), .Q(l8[14]), .QN());
   DFF_X1 \l8_reg[13]  (.D(n_68), .CK(n_3), .Q(l8[13]), .QN());
   DFF_X1 \l8_reg[12]  (.D(n_67), .CK(n_3), .Q(l8[12]), .QN());
   DFF_X1 \l8_reg[11]  (.D(n_66), .CK(n_3), .Q(l8[11]), .QN());
   DFF_X1 \l8_reg[10]  (.D(n_65), .CK(n_3), .Q(l8[10]), .QN());
   DFF_X1 \l8_reg[9]  (.D(n_64), .CK(n_3), .Q(l8[9]), .QN());
   DFF_X1 \l8_reg[8]  (.D(n_63), .CK(n_3), .Q(l8[8]), .QN());
   DFF_X1 \l8_reg[7]  (.D(n_62), .CK(n_3), .Q(l8[7]), .QN());
   DFF_X1 \l8_reg[6]  (.D(n_61), .CK(n_3), .Q(l8[6]), .QN());
   DFF_X1 \l8_reg[5]  (.D(n_60), .CK(n_3), .Q(l8[5]), .QN());
   DFF_X1 \l8_reg[4]  (.D(n_59), .CK(n_3), .Q(l8[4]), .QN());
   DFF_X1 \l8_reg[3]  (.D(n_37), .CK(n_3), .Q(l8[3]), .QN());
   DFF_X1 \l8_reg[2]  (.D(n_36), .CK(n_3), .Q(l8[2]), .QN());
   DFF_X1 \l8_reg[1]  (.D(n_35), .CK(n_3), .Q(l8[1]), .QN());
   DFF_X1 \l8_reg[0]  (.D(n_34), .CK(n_3), .Q(l8[0]), .QN());
   CLKGATETST_X1 clk_gate_f8_reg (.CK(clk), .E(start), .SE(1'b0), .GCK(n_0));
   DFF_X1 \f8_reg[24]  (.D(read2[24]), .CK(n_0), .Q(f8[24]), .QN());
   DFF_X1 \f8_reg[23]  (.D(read2[23]), .CK(n_0), .Q(f8[23]), .QN());
   DFF_X1 \f8_reg[22]  (.D(read[22]), .CK(n_0), .Q(f8[22]), .QN());
   DFF_X1 \f8_reg[21]  (.D(read[21]), .CK(n_0), .Q(f8[21]), .QN());
   DFF_X1 \f8_reg[20]  (.D(read[20]), .CK(n_0), .Q(f8[20]), .QN());
   DFF_X1 \f8_reg[19]  (.D(read[19]), .CK(n_0), .Q(f8[19]), .QN());
   DFF_X1 \f8_reg[18]  (.D(read[18]), .CK(n_0), .Q(f8[18]), .QN());
   DFF_X1 \f8_reg[17]  (.D(read[17]), .CK(n_0), .Q(f8[17]), .QN());
   DFF_X1 \f8_reg[16]  (.D(read[16]), .CK(n_0), .Q(f8[16]), .QN());
   DFF_X1 \f8_reg[15]  (.D(read[15]), .CK(n_0), .Q(f8[15]), .QN());
   DFF_X1 \f8_reg[14]  (.D(read[14]), .CK(n_0), .Q(f8[14]), .QN());
   DFF_X1 \f8_reg[13]  (.D(read[13]), .CK(n_0), .Q(f8[13]), .QN());
   DFF_X1 \f8_reg[12]  (.D(read[12]), .CK(n_0), .Q(f8[12]), .QN());
   DFF_X1 \f8_reg[11]  (.D(read[11]), .CK(n_0), .Q(f8[11]), .QN());
   DFF_X1 \f8_reg[10]  (.D(read[10]), .CK(n_0), .Q(f8[10]), .QN());
   DFF_X1 \f8_reg[9]  (.D(read[9]), .CK(n_0), .Q(f8[9]), .QN());
   DFF_X1 \f8_reg[8]  (.D(read[8]), .CK(n_0), .Q(f8[8]), .QN());
   DFF_X1 \f8_reg[7]  (.D(read[7]), .CK(n_0), .Q(f8[7]), .QN());
   DFF_X1 \f8_reg[6]  (.D(read[6]), .CK(n_0), .Q(f8[6]), .QN());
   DFF_X1 \f8_reg[5]  (.D(read[5]), .CK(n_0), .Q(f8[5]), .QN());
   DFF_X1 \f8_reg[4]  (.D(read[4]), .CK(n_0), .Q(f8[4]), .QN());
   DFF_X1 \f8_reg[3]  (.D(read[3]), .CK(n_0), .Q(f8[3]), .QN());
   DFF_X1 \f8_reg[2]  (.D(read[2]), .CK(n_0), .Q(f8[2]), .QN());
   DFF_X1 \f8_reg[1]  (.D(read[1]), .CK(n_0), .Q(f8[1]), .QN());
   DFF_X1 \f8_reg[0]  (.D(read[0]), .CK(n_0), .Q(f8[0]), .QN());
   DFF_X1 write_en_reg (.D(start), .CK(clk), .Q(write_en), .QN());
   DFF_X1 write_en2_reg (.D(n_88), .CK(clk), .Q(write_en2), .QN());
   DFF_X1 \count_reg[5]  (.D(n_7), .CK(n_3), .Q(count[5]), .QN());
   DFF_X1 \count_reg[4]  (.D(n_6), .CK(n_3), .Q(count[4]), .QN());
   DFF_X1 \count_reg[3]  (.D(n_5), .CK(n_3), .Q(count[3]), .QN());
   DFF_X1 \count_reg[2]  (.D(n_4), .CK(n_3), .Q(count[2]), .QN());
   DFF_X1 \count_reg[1]  (.D(n_2), .CK(n_3), .Q(count[1]), .QN());
   DFF_X1 \count_reg[0]  (.D(n_1), .CK(n_3), .Q(count[0]), .QN());
   DFF_X1 q0_reg (.D(n_81), .CK(n_3), .Q(q0), .QN());
   CLKGATETST_X1 clk_gate_A_reg__2 (.CK(clk), .E(n_82), .SE(1'b0), .GCK(n_3));
   NOR2_X1 i_0_0 (.A1(count[0]), .A2(start), .ZN(n_1));
   AOI21_X1 i_0_1 (.A(n_0_0), .B1(count[0]), .B2(count[1]), .ZN(n_2));
   OAI21_X1 i_0_2 (.A(n_83), .B1(count[0]), .B2(count[1]), .ZN(n_0_0));
   NOR3_X1 i_0_3 (.A1(start), .A2(n_0_6), .A3(n_0_1), .ZN(n_4));
   AOI21_X1 i_0_4 (.A(count[2]), .B1(count[1]), .B2(count[0]), .ZN(n_0_1));
   AOI21_X1 i_0_5 (.A(n_0_2), .B1(n_0_6), .B2(count[3]), .ZN(n_5));
   OAI21_X1 i_0_6 (.A(n_83), .B1(n_0_6), .B2(count[3]), .ZN(n_0_2));
   NOR3_X1 i_0_7 (.A1(start), .A2(n_0_5), .A3(n_0_3), .ZN(n_6));
   AOI21_X1 i_0_8 (.A(count[4]), .B1(count[3]), .B2(n_0_6), .ZN(n_0_3));
   NOR2_X1 i_0_9 (.A1(start), .A2(n_0_4), .ZN(n_7));
   XNOR2_X1 i_0_10 (.A(count[5]), .B(n_0_5), .ZN(n_0_4));
   AND3_X1 i_0_11 (.A1(count[4]), .A2(count[3]), .A3(n_0_6), .ZN(n_0_5));
   AND3_X1 i_0_12 (.A1(count[2]), .A2(count[1]), .A3(count[0]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(n_83), .A2(n_0_39), .ZN(n_8));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_9));
   AOI222_X1 i_0_15 (.A1(n_0_37), .A2(A[1]), .B1(SubM[1]), .B2(n_0_34), .C1(
      AddM[1]), .C2(n_0_35), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_10));
   AOI222_X1 i_0_17 (.A1(n_0_37), .A2(A[2]), .B1(SubM[2]), .B2(n_0_34), .C1(
      AddM[2]), .C2(n_0_35), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_11));
   AOI222_X1 i_0_19 (.A1(n_0_37), .A2(A[3]), .B1(SubM[3]), .B2(n_0_34), .C1(
      AddM[3]), .C2(n_0_35), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_12));
   AOI222_X1 i_0_21 (.A1(n_0_37), .A2(A[4]), .B1(SubM[4]), .B2(n_0_34), .C1(
      AddM[4]), .C2(n_0_35), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_13));
   AOI222_X1 i_0_23 (.A1(n_0_37), .A2(A[5]), .B1(SubM[5]), .B2(n_0_34), .C1(
      AddM[5]), .C2(n_0_35), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_14));
   AOI222_X1 i_0_25 (.A1(n_0_37), .A2(A[6]), .B1(SubM[6]), .B2(n_0_34), .C1(
      AddM[6]), .C2(n_0_35), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_15));
   AOI222_X1 i_0_27 (.A1(n_0_37), .A2(A[7]), .B1(SubM[7]), .B2(n_0_34), .C1(
      AddM[7]), .C2(n_0_35), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_16));
   AOI222_X1 i_0_29 (.A1(n_0_37), .A2(A[8]), .B1(SubM[8]), .B2(n_0_34), .C1(
      AddM[8]), .C2(n_0_35), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_17));
   AOI222_X1 i_0_31 (.A1(n_0_37), .A2(A[9]), .B1(SubM[9]), .B2(n_0_34), .C1(
      AddM[9]), .C2(n_0_35), .ZN(n_0_15));
   INV_X1 i_0_32 (.A(n_0_16), .ZN(n_18));
   AOI222_X1 i_0_33 (.A1(n_0_37), .A2(A[10]), .B1(SubM[10]), .B2(n_0_34), 
      .C1(AddM[10]), .C2(n_0_35), .ZN(n_0_16));
   INV_X1 i_0_34 (.A(n_0_17), .ZN(n_19));
   AOI222_X1 i_0_35 (.A1(n_0_37), .A2(A[11]), .B1(SubM[11]), .B2(n_0_34), 
      .C1(AddM[11]), .C2(n_0_35), .ZN(n_0_17));
   INV_X1 i_0_36 (.A(n_0_18), .ZN(n_20));
   AOI222_X1 i_0_37 (.A1(n_0_37), .A2(A[12]), .B1(SubM[12]), .B2(n_0_34), 
      .C1(AddM[12]), .C2(n_0_35), .ZN(n_0_18));
   INV_X1 i_0_38 (.A(n_0_19), .ZN(n_21));
   AOI222_X1 i_0_39 (.A1(n_0_37), .A2(A[13]), .B1(SubM[13]), .B2(n_0_34), 
      .C1(AddM[13]), .C2(n_0_35), .ZN(n_0_19));
   INV_X1 i_0_40 (.A(n_0_20), .ZN(n_22));
   AOI222_X1 i_0_41 (.A1(n_0_37), .A2(A[14]), .B1(SubM[14]), .B2(n_0_34), 
      .C1(AddM[14]), .C2(n_0_35), .ZN(n_0_20));
   INV_X1 i_0_42 (.A(n_0_21), .ZN(n_23));
   AOI222_X1 i_0_43 (.A1(n_0_37), .A2(A[15]), .B1(SubM[15]), .B2(n_0_34), 
      .C1(AddM[15]), .C2(n_0_35), .ZN(n_0_21));
   INV_X1 i_0_44 (.A(n_0_22), .ZN(n_24));
   AOI222_X1 i_0_45 (.A1(n_0_37), .A2(A[16]), .B1(SubM[16]), .B2(n_0_34), 
      .C1(AddM[16]), .C2(n_0_35), .ZN(n_0_22));
   INV_X1 i_0_46 (.A(n_0_23), .ZN(n_25));
   AOI222_X1 i_0_47 (.A1(n_0_37), .A2(A[17]), .B1(SubM[17]), .B2(n_0_34), 
      .C1(AddM[17]), .C2(n_0_35), .ZN(n_0_23));
   INV_X1 i_0_48 (.A(n_0_24), .ZN(n_26));
   AOI222_X1 i_0_49 (.A1(n_0_37), .A2(A[18]), .B1(SubM[18]), .B2(n_0_34), 
      .C1(AddM[18]), .C2(n_0_35), .ZN(n_0_24));
   INV_X1 i_0_50 (.A(n_0_25), .ZN(n_27));
   AOI222_X1 i_0_51 (.A1(n_0_37), .A2(A[19]), .B1(SubM[19]), .B2(n_0_34), 
      .C1(AddM[19]), .C2(n_0_35), .ZN(n_0_25));
   INV_X1 i_0_52 (.A(n_0_26), .ZN(n_28));
   AOI222_X1 i_0_53 (.A1(n_0_37), .A2(A[20]), .B1(SubM[20]), .B2(n_0_34), 
      .C1(AddM[20]), .C2(n_0_35), .ZN(n_0_26));
   INV_X1 i_0_54 (.A(n_0_27), .ZN(n_29));
   AOI222_X1 i_0_55 (.A1(n_0_37), .A2(A[21]), .B1(SubM[21]), .B2(n_0_34), 
      .C1(AddM[21]), .C2(n_0_35), .ZN(n_0_27));
   INV_X1 i_0_56 (.A(n_0_28), .ZN(n_30));
   AOI222_X1 i_0_57 (.A1(n_0_37), .A2(A[22]), .B1(SubM[22]), .B2(n_0_34), 
      .C1(AddM[22]), .C2(n_0_35), .ZN(n_0_28));
   INV_X1 i_0_58 (.A(n_0_29), .ZN(n_31));
   AOI222_X1 i_0_59 (.A1(n_0_37), .A2(A[23]), .B1(SubM[23]), .B2(n_0_34), 
      .C1(AddM[23]), .C2(n_0_35), .ZN(n_0_29));
   NAND2_X1 i_0_60 (.A1(n_0_30), .A2(n_0_31), .ZN(n_32));
   NAND2_X1 i_0_61 (.A1(n_0_37), .A2(A[24]), .ZN(n_0_30));
   INV_X1 i_0_62 (.A(n_0_31), .ZN(n_33));
   AOI22_X1 i_0_63 (.A1(AddM[24]), .A2(n_0_35), .B1(n_0_34), .B2(SubM[24]), 
      .ZN(n_0_31));
   MUX2_X1 i_0_64 (.A(l8[1]), .B(read2[0]), .S(start), .Z(n_34));
   MUX2_X1 i_0_65 (.A(l8[2]), .B(read2[1]), .S(start), .Z(n_35));
   MUX2_X1 i_0_66 (.A(l8[3]), .B(read2[2]), .S(start), .Z(n_36));
   MUX2_X1 i_0_67 (.A(l8[4]), .B(read2[3]), .S(start), .Z(n_37));
   MUX2_X1 i_0_68 (.A(l8[5]), .B(read2[4]), .S(start), .Z(n_59));
   MUX2_X1 i_0_69 (.A(l8[6]), .B(read2[5]), .S(start), .Z(n_60));
   MUX2_X1 i_0_70 (.A(l8[7]), .B(read2[6]), .S(start), .Z(n_61));
   MUX2_X1 i_0_71 (.A(l8[8]), .B(read2[7]), .S(start), .Z(n_62));
   MUX2_X1 i_0_72 (.A(l8[9]), .B(read2[8]), .S(start), .Z(n_63));
   MUX2_X1 i_0_73 (.A(l8[10]), .B(read2[9]), .S(start), .Z(n_64));
   MUX2_X1 i_0_74 (.A(l8[11]), .B(read2[10]), .S(start), .Z(n_65));
   MUX2_X1 i_0_75 (.A(l8[12]), .B(read2[11]), .S(start), .Z(n_66));
   MUX2_X1 i_0_76 (.A(l8[13]), .B(read2[12]), .S(start), .Z(n_67));
   MUX2_X1 i_0_77 (.A(l8[14]), .B(read2[13]), .S(start), .Z(n_68));
   MUX2_X1 i_0_78 (.A(l8[15]), .B(read2[14]), .S(start), .Z(n_69));
   MUX2_X1 i_0_79 (.A(l8[16]), .B(read2[15]), .S(start), .Z(n_70));
   MUX2_X1 i_0_80 (.A(l8[17]), .B(read2[16]), .S(start), .Z(n_71));
   MUX2_X1 i_0_81 (.A(l8[18]), .B(read2[17]), .S(start), .Z(n_72));
   MUX2_X1 i_0_82 (.A(l8[19]), .B(read2[18]), .S(start), .Z(n_73));
   MUX2_X1 i_0_83 (.A(l8[20]), .B(read2[19]), .S(start), .Z(n_74));
   MUX2_X1 i_0_84 (.A(l8[21]), .B(read2[20]), .S(start), .Z(n_75));
   MUX2_X1 i_0_85 (.A(l8[22]), .B(read2[21]), .S(start), .Z(n_76));
   MUX2_X1 i_0_86 (.A(l8[23]), .B(read2[22]), .S(start), .Z(n_77));
   MUX2_X1 i_0_87 (.A(l8[24]), .B(read2[23]), .S(start), .Z(n_78));
   NAND2_X1 i_0_88 (.A1(n_0_33), .A2(n_0_32), .ZN(n_79));
   AOI22_X1 i_0_89 (.A1(AddM[0]), .A2(n_0_35), .B1(n_0_34), .B2(SubM[0]), 
      .ZN(n_0_32));
   AOI22_X1 i_0_90 (.A1(n_0_37), .A2(A[0]), .B1(start), .B2(read2[24]), .ZN(
      n_0_33));
   NOR3_X1 i_0_91 (.A1(n_0_42), .A2(start), .A3(q0), .ZN(n_0_34));
   AND3_X1 i_0_92 (.A1(n_0_42), .A2(n_83), .A3(q0), .ZN(n_0_35));
   NAND2_X1 i_0_93 (.A1(n_83), .A2(n_0_36), .ZN(n_80));
   NAND2_X1 i_0_94 (.A1(n_0_39), .A2(n_0_38), .ZN(n_0_36));
   NOR2_X1 i_0_95 (.A1(n_0_38), .A2(start), .ZN(n_0_37));
   XNOR2_X1 i_0_96 (.A(q0), .B(n_0_42), .ZN(n_0_38));
   NOR2_X1 i_0_97 (.A1(n_0_42), .A2(start), .ZN(n_81));
   OR2_X1 i_0_98 (.A1(n_0_39), .A2(start), .ZN(n_82));
   NAND3_X1 i_0_99 (.A1(count[4]), .A2(count[3]), .A3(n_0_40), .ZN(n_0_39));
   NOR4_X1 i_0_100 (.A1(count[2]), .A2(n_0_41), .A3(count[1]), .A4(count[5]), 
      .ZN(n_0_40));
   INV_X1 i_0_101 (.A(start), .ZN(n_83));
   INV_X1 i_0_102 (.A(count[0]), .ZN(n_0_41));
   INV_X1 i_0_103 (.A(l8[0]), .ZN(n_0_42));
   MUX2_X1 \A_reg[24]_enable_mux_0  (.A(A[24]), .B(n_33), .S(n_80), .Z(n_87));
   MUX2_X1 write_en2_reg_enable_mux_0 (.A(write_en2), .B(n_83), .S(n_8), 
      .Z(n_88));
   datapath__0_24 i_17 (.f8(f8), .p_0({n_86, n_85, n_84, n_58, n_57, n_56, n_55, 
      n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, uc_56}));
endmodule

module normalize(mantissa, mantissaOutFinal, carry);
   input [47:0]mantissa;
   output [22:0]mantissaOutFinal;
   output carry;

   INV_X1 i_0_0 (.A(mantissa[46]), .ZN(carry));
   MUX2_X1 i_0_1 (.A(mantissa[24]), .B(mantissa[23]), .S(mantissa[46]), .Z(
      mantissaOutFinal[0]));
   MUX2_X1 i_0_2 (.A(mantissa[25]), .B(mantissa[24]), .S(mantissa[46]), .Z(
      mantissaOutFinal[1]));
   MUX2_X1 i_0_3 (.A(mantissa[26]), .B(mantissa[25]), .S(mantissa[46]), .Z(
      mantissaOutFinal[2]));
   MUX2_X1 i_0_4 (.A(mantissa[27]), .B(mantissa[26]), .S(mantissa[46]), .Z(
      mantissaOutFinal[3]));
   MUX2_X1 i_0_5 (.A(mantissa[28]), .B(mantissa[27]), .S(mantissa[46]), .Z(
      mantissaOutFinal[4]));
   MUX2_X1 i_0_6 (.A(mantissa[29]), .B(mantissa[28]), .S(mantissa[46]), .Z(
      mantissaOutFinal[5]));
   MUX2_X1 i_0_7 (.A(mantissa[30]), .B(mantissa[29]), .S(mantissa[46]), .Z(
      mantissaOutFinal[6]));
   MUX2_X1 i_0_8 (.A(mantissa[31]), .B(mantissa[30]), .S(mantissa[46]), .Z(
      mantissaOutFinal[7]));
   MUX2_X1 i_0_9 (.A(mantissa[32]), .B(mantissa[31]), .S(mantissa[46]), .Z(
      mantissaOutFinal[8]));
   MUX2_X1 i_0_10 (.A(mantissa[33]), .B(mantissa[32]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[9]));
   MUX2_X1 i_0_11 (.A(mantissa[34]), .B(mantissa[33]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[10]));
   MUX2_X1 i_0_12 (.A(mantissa[35]), .B(mantissa[34]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[11]));
   MUX2_X1 i_0_13 (.A(mantissa[36]), .B(mantissa[35]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[12]));
   MUX2_X1 i_0_14 (.A(mantissa[37]), .B(mantissa[36]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[13]));
   MUX2_X1 i_0_15 (.A(mantissa[38]), .B(mantissa[37]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[14]));
   MUX2_X1 i_0_16 (.A(mantissa[39]), .B(mantissa[38]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[15]));
   MUX2_X1 i_0_17 (.A(mantissa[40]), .B(mantissa[39]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[16]));
   MUX2_X1 i_0_18 (.A(mantissa[41]), .B(mantissa[40]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[17]));
   MUX2_X1 i_0_19 (.A(mantissa[42]), .B(mantissa[41]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[18]));
   MUX2_X1 i_0_20 (.A(mantissa[43]), .B(mantissa[42]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[19]));
   MUX2_X1 i_0_21 (.A(mantissa[44]), .B(mantissa[43]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[20]));
   MUX2_X1 i_0_22 (.A(mantissa[45]), .B(mantissa[44]), .S(mantissa[46]), 
      .Z(mantissaOutFinal[21]));
   AND2_X1 i_0_23 (.A1(mantissa[45]), .A2(mantissa[46]), .ZN(
      mantissaOutFinal[22]));
endmodule

module full_adder__0_32(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
   AND2_X1 i_0_1 (.A1(i_bit2), .A2(i_bit1), .ZN(o_carry));
endmodule

module full_adder__0_36(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_40(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_44(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_48(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_52(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_56(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(i_carry), .Z(o_sum));
endmodule

module ripple_adder(i_add1, i_add2, o_result, o_carry);
   input [7:0]i_add1;
   input [7:0]i_add2;
   output [7:0]o_result;
   output o_carry;

   full_adder__0_32 genblk1_0_full_adder_inst (.i_bit1(i_add1[0]), .i_bit2(
      i_add2[0]), .i_carry(), .o_sum(o_result[0]), .o_carry(n_0));
   full_adder__0_36 genblk1_1_full_adder_inst (.i_bit1(i_add1[1]), .i_bit2(
      i_add2[1]), .i_carry(n_0), .o_sum(o_result[1]), .o_carry(n_1));
   full_adder__0_40 genblk1_2_full_adder_inst (.i_bit1(i_add1[2]), .i_bit2(
      i_add2[2]), .i_carry(n_1), .o_sum(o_result[2]), .o_carry(n_2));
   full_adder__0_44 genblk1_3_full_adder_inst (.i_bit1(i_add1[3]), .i_bit2(
      i_add2[3]), .i_carry(n_2), .o_sum(o_result[3]), .o_carry(n_3));
   full_adder__0_48 genblk1_4_full_adder_inst (.i_bit1(i_add1[4]), .i_bit2(
      i_add2[4]), .i_carry(n_3), .o_sum(o_result[4]), .o_carry(n_4));
   full_adder__0_52 genblk1_5_full_adder_inst (.i_bit1(i_add1[5]), .i_bit2(
      i_add2[5]), .i_carry(n_4), .o_sum(o_result[5]), .o_carry(n_5));
   full_adder__0_56 genblk1_6_full_adder_inst (.i_bit1(i_add1[6]), .i_bit2(
      i_add2[6]), .i_carry(n_5), .o_sum(o_result[6]), .o_carry(n_6));
   full_adder genblk1_7_full_adder_inst (.i_bit1(i_add1[7]), .i_bit2(i_add2[7]), 
      .i_carry(n_6), .o_sum(o_result[7]), .o_carry());
endmodule

module fp_multiplier(inputA, inputB, leading1, bias, result, over_flow, 
      under_flow, clk, start, left_bias);
   input [31:0]inputA;
   input [31:0]inputB;
   input [1:0]leading1;
   input [7:0]bias;
   output [31:0]result;
   output over_flow;
   output under_flow;
   input clk;
   input start;
   input [6:0]left_bias;

   wire [31:0]no_result;
   wire control_signal;
   wire finalSign;
   wire [7:0]addition_exp;
   wire n_0_32;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_23;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire carry_normalize;
   wire [22:0]mantissa_out;
   wire [7:0]output_exp;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;

   assign under_flow = 1'b0;

   subnormal subnormal_inst (.inputA({inputA[30], inputA[29], inputA[28], 
      inputA[27], inputA[26], inputA[25], inputA[24], inputA[23]}), .inputB({
      inputB[30], inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], 
      inputB[24], inputB[23]}), .overflow(control_signal), .signal(), .result(
      no_result));
   xor_module xor_inst (.sign1(inputA[31]), .sign2(inputB[31]), .sign_out(
      finalSign));
   ripple_adder__0_89 adder_inst1 (.i_add1({inputA[30], inputA[29], inputA[28], 
      inputA[27], inputA[26], inputA[25], inputA[24], inputA[23]}), .i_add2({
      inputB[30], inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], 
      inputB[24], inputB[23]}), .o_result(addition_exp), .o_carry());
   ripple_adder__0_122 adder_inst2 (.i_add1(addition_exp), .i_add2(bias), 
      .o_result({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24}), 
      .o_carry(n_0_32));
   BoothAlgo multiplier_inst (.M({leading1[1], leading1[0], inputA[22], 
      inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
      inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], 
      inputA[9], inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], 
      inputA[3], inputA[2], inputA[1], inputA[0]}), .Q({uc_0, uc_1, inputB[22], 
      inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
      inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], 
      inputB[9], inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], 
      inputB[3], inputB[2], inputB[1], inputB[0]}), .result({uc_2, uc_3, uc_4, 
      n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
      n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
      n_0_3, n_0_2, n_0_1, n_0_0, n_0_23, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, 
      uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, 
      uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27}), .clk(clk), .start(start));
   normalize normalizer_inst (.mantissa({uc_28, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
      n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, 
      n_0_23, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, 
      uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, 
      uc_48, uc_49, uc_50, uc_51}), .mantissaOutFinal(mantissa_out), .carry(
      carry_normalize));
   ripple_adder adder_inst3 (.i_add1({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24}), .i_add2({left_bias[6], left_bias[5], 
      left_bias[4], left_bias[3], left_bias[2], left_bias[1], left_bias[0], 
      carry_normalize}), .o_result(output_exp), .o_carry());
   OAI21_X1 i_0_0_0 (.A(n_0_0_0), .B1(n_0_0_1), .B2(n_0_0_2), .ZN(over_flow));
   NOR2_X1 i_0_0_1 (.A1(control_signal), .A2(n_0_32), .ZN(n_0_0_0));
   NAND4_X1 i_0_0_2 (.A1(output_exp[7]), .A2(output_exp[6]), .A3(output_exp[5]), 
      .A4(output_exp[4]), .ZN(n_0_0_1));
   NAND4_X1 i_0_0_3 (.A1(output_exp[3]), .A2(output_exp[2]), .A3(output_exp[1]), 
      .A4(output_exp[0]), .ZN(n_0_0_2));
   MUX2_X1 i_0_0_4 (.A(mantissa_out[0]), .B(no_result[0]), .S(control_signal), 
      .Z(result[0]));
   MUX2_X1 i_0_0_5 (.A(mantissa_out[1]), .B(no_result[1]), .S(control_signal), 
      .Z(result[1]));
   MUX2_X1 i_0_0_6 (.A(mantissa_out[2]), .B(no_result[2]), .S(control_signal), 
      .Z(result[2]));
   MUX2_X1 i_0_0_7 (.A(mantissa_out[3]), .B(no_result[3]), .S(control_signal), 
      .Z(result[3]));
   MUX2_X1 i_0_0_8 (.A(mantissa_out[4]), .B(no_result[4]), .S(control_signal), 
      .Z(result[4]));
   MUX2_X1 i_0_0_9 (.A(mantissa_out[5]), .B(no_result[5]), .S(control_signal), 
      .Z(result[5]));
   MUX2_X1 i_0_0_10 (.A(mantissa_out[6]), .B(no_result[6]), .S(control_signal), 
      .Z(result[6]));
   MUX2_X1 i_0_0_11 (.A(mantissa_out[7]), .B(no_result[7]), .S(control_signal), 
      .Z(result[7]));
   MUX2_X1 i_0_0_12 (.A(mantissa_out[8]), .B(no_result[8]), .S(control_signal), 
      .Z(result[8]));
   MUX2_X1 i_0_0_13 (.A(mantissa_out[9]), .B(no_result[9]), .S(control_signal), 
      .Z(result[9]));
   MUX2_X1 i_0_0_14 (.A(mantissa_out[10]), .B(no_result[10]), .S(control_signal), 
      .Z(result[10]));
   MUX2_X1 i_0_0_15 (.A(mantissa_out[11]), .B(no_result[11]), .S(control_signal), 
      .Z(result[11]));
   MUX2_X1 i_0_0_16 (.A(mantissa_out[12]), .B(no_result[12]), .S(control_signal), 
      .Z(result[12]));
   MUX2_X1 i_0_0_17 (.A(mantissa_out[13]), .B(no_result[13]), .S(control_signal), 
      .Z(result[13]));
   MUX2_X1 i_0_0_18 (.A(mantissa_out[14]), .B(no_result[14]), .S(control_signal), 
      .Z(result[14]));
   MUX2_X1 i_0_0_19 (.A(mantissa_out[15]), .B(no_result[15]), .S(control_signal), 
      .Z(result[15]));
   MUX2_X1 i_0_0_20 (.A(mantissa_out[16]), .B(no_result[16]), .S(control_signal), 
      .Z(result[16]));
   MUX2_X1 i_0_0_21 (.A(mantissa_out[17]), .B(no_result[17]), .S(control_signal), 
      .Z(result[17]));
   MUX2_X1 i_0_0_22 (.A(mantissa_out[18]), .B(no_result[18]), .S(control_signal), 
      .Z(result[18]));
   MUX2_X1 i_0_0_23 (.A(mantissa_out[19]), .B(no_result[19]), .S(control_signal), 
      .Z(result[19]));
   MUX2_X1 i_0_0_24 (.A(mantissa_out[20]), .B(no_result[20]), .S(control_signal), 
      .Z(result[20]));
   MUX2_X1 i_0_0_25 (.A(mantissa_out[21]), .B(no_result[21]), .S(control_signal), 
      .Z(result[21]));
   MUX2_X1 i_0_0_26 (.A(mantissa_out[22]), .B(no_result[22]), .S(control_signal), 
      .Z(result[22]));
   MUX2_X1 i_0_0_27 (.A(output_exp[0]), .B(no_result[23]), .S(control_signal), 
      .Z(result[23]));
   MUX2_X1 i_0_0_28 (.A(output_exp[1]), .B(no_result[24]), .S(control_signal), 
      .Z(result[24]));
   MUX2_X1 i_0_0_29 (.A(output_exp[2]), .B(no_result[25]), .S(control_signal), 
      .Z(result[25]));
   MUX2_X1 i_0_0_30 (.A(output_exp[3]), .B(no_result[26]), .S(control_signal), 
      .Z(result[26]));
   MUX2_X1 i_0_0_31 (.A(output_exp[4]), .B(no_result[27]), .S(control_signal), 
      .Z(result[27]));
   MUX2_X1 i_0_0_32 (.A(output_exp[5]), .B(no_result[28]), .S(control_signal), 
      .Z(result[28]));
   MUX2_X1 i_0_0_33 (.A(output_exp[6]), .B(no_result[29]), .S(control_signal), 
      .Z(result[29]));
   MUX2_X1 i_0_0_34 (.A(output_exp[7]), .B(no_result[30]), .S(control_signal), 
      .Z(result[30]));
   MUX2_X1 i_0_0_35 (.A(finalSign), .B(no_result[31]), .S(control_signal), 
      .Z(result[31]));
endmodule
